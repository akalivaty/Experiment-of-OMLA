//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1059, new_n1060;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  NAND3_X1  g002(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G183gat), .B2(G190gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206));
  AND2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(KEYINPUT24), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n203), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n205), .A2(new_n209), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(new_n203), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n215), .A2(new_n221), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(KEYINPUT23), .B2(new_n212), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n218), .A2(new_n220), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT66), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(new_n215), .A3(new_n231), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n237), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT28), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n245), .B2(G190gat), .ZN(new_n246));
  INV_X1    g045(.A(G190gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(KEYINPUT28), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n227), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n237), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT67), .B1(new_n236), .B2(new_n237), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n227), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n226), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G113gat), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G120gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT1), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G127gat), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G127gat), .A2(G134gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT69), .B1(new_n264), .B2(new_n265), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n256), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n259), .A2(G120gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n257), .A2(G113gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n273), .B1(new_n276), .B2(new_n266), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n261), .B2(new_n274), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n269), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n255), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n226), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n284), .B2(new_n253), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n279), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G227gat), .ZN(new_n288));
  INV_X1    g087(.A(G233gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT34), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT71), .B1(new_n287), .B2(new_n290), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298));
  INV_X1    g097(.A(new_n290), .ZN(new_n299));
  AOI211_X1 g098(.A(new_n298), .B(new_n299), .C1(new_n281), .C2(new_n286), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT32), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT33), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n297), .B2(new_n300), .ZN(new_n303));
  XOR2_X1   g102(.A(G15gat), .B(G43gat), .Z(new_n304));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n253), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n279), .B1(new_n309), .B2(new_n226), .ZN(new_n310));
  AOI211_X1 g109(.A(new_n280), .B(new_n282), .C1(new_n284), .C2(new_n253), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n290), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n298), .ZN(new_n313));
  OAI211_X1 g112(.A(KEYINPUT71), .B(new_n290), .C1(new_n310), .C2(new_n311), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT33), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  INV_X1    g115(.A(new_n306), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n296), .B1(new_n307), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  INV_X1    g119(.A(new_n296), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n322));
  AOI221_X4 g121(.A(new_n308), .B1(KEYINPUT33), .B2(new_n306), .C1(new_n313), .C2(new_n314), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n318), .A3(new_n296), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G141gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n332), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n334), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT77), .B(G148gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(G141gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n331), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n338), .B2(new_n329), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT78), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n335), .A2(KEYINPUT77), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G148gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n334), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n331), .B1(new_n330), .B2(KEYINPUT2), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n340), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT78), .B1(new_n343), .B2(new_n345), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n347), .A3(new_n353), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n339), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT79), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365));
  AND2_X1   g164(.A1(G211gat), .A2(G218gat), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n364), .A2(new_n365), .B1(new_n366), .B2(KEYINPUT22), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n368));
  NOR2_X1   g167(.A1(G211gat), .A2(G218gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n366), .A2(new_n369), .ZN(new_n371));
  INV_X1    g170(.A(G197gat), .ZN(new_n372));
  INV_X1    g171(.A(G204gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT22), .ZN(new_n375));
  NAND2_X1  g174(.A1(G211gat), .A2(G218gat), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n374), .A2(new_n363), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n371), .B1(new_n377), .B2(KEYINPUT74), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n362), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n361), .A3(new_n380), .ZN(new_n381));
  AOI211_X1 g180(.A(KEYINPUT3), .B(new_n339), .C1(new_n358), .C2(new_n359), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n379), .B1(new_n382), .B2(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n379), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n362), .B(new_n340), .C1(new_n346), .C2(new_n354), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  INV_X1    g190(.A(G218gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT80), .B1(new_n393), .B2(new_n376), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n367), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n366), .B2(new_n369), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n371), .A2(KEYINPUT80), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n389), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n360), .B1(new_n402), .B2(new_n362), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n384), .B1(new_n390), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n406), .B(new_n384), .C1(new_n390), .C2(new_n403), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n386), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n409));
  OAI21_X1  g208(.A(G22gat), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI211_X1 g209(.A(KEYINPUT82), .B(new_n386), .C1(new_n405), .C2(new_n407), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n328), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G78gat), .B(G106gat), .Z(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT31), .B(G50gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n417));
  INV_X1    g216(.A(new_n407), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n395), .A2(new_n398), .B1(KEYINPUT80), .B2(new_n371), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n362), .B1(new_n419), .B2(KEYINPUT29), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n355), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n360), .B2(new_n362), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n387), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n406), .B1(new_n423), .B2(new_n384), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n408), .A2(KEYINPUT84), .A3(new_n416), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n415), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n417), .B1(new_n418), .B2(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT82), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n409), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT83), .A4(G22gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n412), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n408), .A2(new_n416), .ZN(new_n435));
  INV_X1    g234(.A(new_n425), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n415), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n320), .A2(new_n327), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n283), .A2(new_n443), .A3(new_n226), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(KEYINPUT29), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n444), .B(new_n379), .C1(new_n285), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n283), .A2(new_n226), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n285), .A2(new_n443), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n447), .B(KEYINPUT75), .C1(new_n449), .C2(new_n379), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n285), .A2(new_n443), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n387), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n450), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n450), .B2(new_n455), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n450), .A2(new_n455), .ZN(new_n465));
  AND4_X1   g264(.A1(KEYINPUT76), .A2(new_n465), .A3(KEYINPUT30), .A4(new_n458), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT76), .B1(new_n461), .B2(KEYINPUT30), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT4), .B1(new_n360), .B2(new_n279), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n279), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n357), .A2(new_n361), .A3(KEYINPUT3), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n382), .A2(new_n279), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g273(.A1(G225gat), .A2(G233gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n357), .A2(new_n361), .A3(new_n280), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n360), .A2(new_n279), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n475), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n471), .A2(new_n472), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n470), .A2(new_n469), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n475), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G1gat), .B(G29gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT0), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G85gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n485), .A3(new_n490), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n491), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n468), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n202), .B1(new_n442), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n439), .A2(new_n441), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n307), .A2(new_n318), .A3(new_n296), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT91), .B(KEYINPUT35), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n501), .A2(new_n319), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n500), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n434), .A2(new_n440), .A3(new_n437), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n440), .B1(new_n434), .B2(new_n437), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n498), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n451), .A2(new_n379), .A3(new_n452), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT89), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n449), .A2(new_n513), .A3(new_n379), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n444), .B1(new_n285), .B2(new_n446), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n387), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT38), .B1(new_n517), .B2(KEYINPUT37), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n465), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n459), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n497), .A2(new_n510), .A3(new_n462), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n495), .A2(new_n496), .A3(new_n462), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n518), .A2(new_n459), .A3(new_n520), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT90), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n459), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n465), .A2(new_n519), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT38), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n522), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n477), .A2(new_n475), .A3(new_n478), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n530), .A2(KEYINPUT88), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT39), .B1(new_n530), .B2(KEYINPUT88), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n482), .A2(new_n483), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT86), .A3(new_n480), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT86), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n473), .B2(new_n475), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT86), .B1(new_n534), .B2(new_n480), .ZN(new_n540));
  AOI211_X1 g339(.A(new_n536), .B(new_n475), .C1(new_n482), .C2(new_n483), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n538), .A2(new_n542), .A3(KEYINPUT40), .A4(new_n490), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n538), .A2(new_n490), .A3(new_n542), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT40), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n544), .A2(new_n545), .B1(new_n491), .B2(new_n486), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n468), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n505), .B2(new_n506), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n509), .B1(new_n529), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n327), .B2(new_n320), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT36), .B1(new_n324), .B2(new_n326), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n499), .A2(new_n504), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT105), .ZN(new_n556));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT101), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT41), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  OR2_X1    g360(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(G85gat), .A3(G92gat), .A4(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n565));
  NOR2_X1   g364(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  OAI22_X1  g367(.A1(new_n565), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G99gat), .ZN(new_n571));
  INV_X1    g370(.A(G106gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT8), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT103), .B(G92gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(G85gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n561), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT8), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(G99gat), .B2(G106gat), .ZN(new_n578));
  AND2_X1   g377(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(KEYINPUT103), .A2(G92gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n581), .B2(new_n567), .ZN(new_n582));
  INV_X1    g381(.A(new_n561), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n564), .A4(new_n569), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT104), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n576), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(KEYINPUT104), .B(new_n561), .C1(new_n570), .C2(new_n575), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT14), .ZN(new_n589));
  INV_X1    g388(.A(G29gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n592));
  AOI21_X1  g391(.A(G36gat), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT15), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G36gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n592), .ZN(new_n598));
  NOR2_X1   g397(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT15), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n594), .ZN(new_n602));
  XNOR2_X1  g401(.A(G43gat), .B(G50gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n605), .B(KEYINPUT15), .C1(new_n593), .C2(new_n595), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n560), .B1(new_n588), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n604), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n604), .B2(new_n606), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n587), .B(new_n586), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n556), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT106), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n558), .A2(new_n559), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n263), .ZN(new_n617));
  INV_X1    g416(.A(G162gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT107), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n608), .A2(new_n612), .A3(new_n556), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n613), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT107), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n624), .B(new_n619), .C1(new_n613), .C2(new_n614), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n615), .B2(new_n619), .ZN(new_n627));
  INV_X1    g426(.A(new_n625), .ZN(new_n628));
  OAI22_X1  g427(.A1(new_n627), .A2(new_n628), .B1(new_n613), .B2(new_n622), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n416), .A2(G15gat), .ZN(new_n632));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(G22gat), .ZN(new_n634));
  INV_X1    g433(.A(G1gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT16), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G8gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G15gat), .B(G22gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(G1gat), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n631), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(G8gat), .B1(new_n640), .B2(new_n636), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n632), .A2(new_n634), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n635), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(KEYINPUT93), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(KEYINPUT92), .A3(new_n637), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT92), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n634), .A3(new_n636), .A4(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(G8gat), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n642), .A2(new_n646), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT21), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(G57gat), .ZN(new_n655));
  INV_X1    g454(.A(G64gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G71gat), .B(G78gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G71gat), .ZN(new_n660));
  INV_X1    g459(.A(G78gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(KEYINPUT9), .ZN(new_n662));
  NAND2_X1  g461(.A1(G71gat), .A2(G78gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n655), .A2(KEYINPUT98), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(G64gat), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n655), .A2(KEYINPUT97), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n656), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n659), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n651), .B1(new_n652), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n652), .ZN(new_n674));
  XNOR2_X1  g473(.A(G127gat), .B(G155gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n673), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G231gat), .A2(G233gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT99), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G183gat), .B(G211gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n677), .B(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT108), .B1(new_n630), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n684), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(new_n629), .A3(new_n687), .A4(new_n626), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n610), .A2(new_n611), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n604), .A2(new_n606), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT94), .B1(new_n691), .B2(new_n651), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n647), .A2(new_n650), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n639), .A2(new_n641), .A3(new_n631), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT93), .B1(new_n643), .B2(new_n645), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT94), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n607), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n690), .A2(new_n651), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(G229gat), .A2(G233gat), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n699), .A2(KEYINPUT95), .A3(KEYINPUT18), .A4(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT95), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n651), .B1(new_n610), .B2(new_n611), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n691), .A2(new_n651), .A3(KEYINPUT94), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n697), .B1(new_n696), .B2(new_n607), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n703), .B(new_n700), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT18), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n707), .ZN(new_n710));
  OAI22_X1  g509(.A1(new_n704), .A2(new_n705), .B1(new_n696), .B2(new_n607), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n700), .B(KEYINPUT13), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(G113gat), .B(G141gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G197gat), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT11), .B(G169gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT12), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT96), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n709), .A2(new_n714), .A3(new_n722), .A4(new_n719), .ZN(new_n723));
  INV_X1    g522(.A(new_n719), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n714), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n721), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n586), .A2(new_n671), .A3(new_n587), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT10), .ZN(new_n728));
  INV_X1    g527(.A(new_n671), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n576), .A3(new_n584), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n727), .A2(KEYINPUT109), .A3(new_n730), .A4(new_n728), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(KEYINPUT10), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n588), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(G230gat), .A2(G233gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n727), .A2(new_n730), .ZN(new_n742));
  INV_X1    g541(.A(new_n740), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(G120gat), .B(G148gat), .Z(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT110), .ZN(new_n746));
  XNOR2_X1  g545(.A(G176gat), .B(G204gat), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n746), .B(new_n747), .Z(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n741), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n733), .A2(new_n734), .B1(new_n588), .B2(new_n737), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n751), .B2(new_n743), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n689), .A2(new_n726), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n554), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n497), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n635), .ZN(G1324gat));
  INV_X1    g558(.A(new_n468), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT16), .B(G8gat), .Z(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n638), .B2(new_n761), .ZN(new_n764));
  MUX2_X1   g563(.A(new_n763), .B(new_n764), .S(KEYINPUT42), .Z(G1325gat));
  NOR3_X1   g564(.A1(new_n501), .A2(new_n319), .A3(KEYINPUT73), .ZN(new_n766));
  INV_X1    g565(.A(new_n320), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT36), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769));
  INV_X1    g568(.A(new_n552), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT111), .B1(new_n551), .B2(new_n552), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G15gat), .B1(new_n756), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n501), .A2(new_n319), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n633), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n756), .B2(new_n776), .ZN(G1326gat));
  NOR2_X1   g576(.A1(new_n756), .A2(new_n500), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT43), .B(G22gat), .Z(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1327gat));
  NAND2_X1  g579(.A1(new_n327), .A2(new_n320), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n500), .A3(new_n498), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT35), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n503), .A2(new_n498), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n500), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n544), .A2(new_n545), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n786), .A2(new_n492), .A3(new_n543), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n439), .A2(new_n441), .B1(new_n787), .B2(new_n468), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n522), .A2(new_n525), .A3(new_n528), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(new_n789), .B1(new_n507), .B2(new_n508), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n768), .A2(new_n770), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n783), .A2(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n630), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n726), .A2(new_n686), .A3(new_n754), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n590), .A3(new_n497), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT45), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT44), .B1(new_n792), .B2(new_n793), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n549), .B1(new_n772), .B2(new_n771), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n782), .A2(KEYINPUT35), .B1(new_n784), .B2(new_n500), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n795), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G29gat), .B1(new_n805), .B2(new_n757), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n798), .A2(new_n806), .ZN(G1328gat));
  NAND3_X1  g606(.A1(new_n796), .A2(new_n597), .A3(new_n468), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT46), .Z(new_n809));
  OAI21_X1  g608(.A(G36gat), .B1(new_n805), .B2(new_n760), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1329gat));
  AOI21_X1  g610(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n551), .A2(KEYINPUT111), .A3(new_n552), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n800), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n773), .A2(new_n790), .ZN(new_n816));
  INV_X1    g615(.A(new_n802), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n554), .B2(new_n630), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n814), .B(new_n794), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n804), .A2(new_n823), .A3(new_n814), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(G43gat), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n796), .ZN(new_n826));
  INV_X1    g625(.A(new_n775), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n826), .A2(G43gat), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT47), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n821), .A2(G43gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n832), .B2(new_n828), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1330gat));
  INV_X1    g633(.A(KEYINPUT48), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n837));
  INV_X1    g636(.A(G50gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n804), .B2(new_n507), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n507), .A2(new_n838), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT113), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n796), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n836), .B(new_n837), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n507), .B(new_n794), .C1(new_n818), .C2(new_n820), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G50gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n846), .A2(KEYINPUT114), .A3(new_n835), .A4(new_n842), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n844), .A2(new_n847), .ZN(G1331gat));
  NAND2_X1  g647(.A1(new_n816), .A2(new_n817), .ZN(new_n849));
  INV_X1    g648(.A(new_n726), .ZN(new_n850));
  INV_X1    g649(.A(new_n754), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n689), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n802), .B1(new_n773), .B2(new_n790), .ZN(new_n855));
  INV_X1    g654(.A(new_n852), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n497), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n667), .A2(G57gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n669), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n860), .B(new_n862), .ZN(G1332gat));
  XNOR2_X1  g662(.A(KEYINPUT49), .B(G64gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n468), .A3(new_n864), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n858), .A2(new_n760), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1333gat));
  OAI21_X1  g666(.A(G71gat), .B1(new_n858), .B2(new_n773), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n857), .A3(new_n660), .A4(new_n775), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(KEYINPUT50), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1334gat));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n500), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(new_n661), .ZN(G1335gat));
  NAND2_X1  g675(.A1(new_n726), .A2(new_n684), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT116), .Z(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n851), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n818), .B2(new_n820), .ZN(new_n880));
  OAI21_X1  g679(.A(G85gat), .B1(new_n880), .B2(new_n757), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n878), .A2(new_n793), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n849), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n849), .A2(KEYINPUT51), .A3(new_n882), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n497), .A2(new_n567), .A3(new_n754), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(G1336gat));
  OAI21_X1  g688(.A(new_n574), .B1(new_n880), .B2(new_n760), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n468), .A2(new_n568), .A3(new_n754), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n890), .B(new_n891), .C1(new_n887), .C2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n885), .B2(new_n886), .ZN(new_n894));
  INV_X1    g693(.A(new_n879), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n799), .B2(new_n803), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n581), .B1(new_n896), .B2(new_n468), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT52), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(G1337gat));
  OAI21_X1  g698(.A(G99gat), .B1(new_n880), .B2(new_n773), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n775), .A2(new_n571), .A3(new_n754), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n887), .B2(new_n901), .ZN(G1338gat));
  OAI21_X1  g701(.A(G106gat), .B1(new_n880), .B2(new_n500), .ZN(new_n903));
  XNOR2_X1  g702(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n507), .A2(new_n572), .A3(new_n754), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n903), .B(new_n904), .C1(new_n887), .C2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n904), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n885), .B2(new_n886), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n572), .B1(new_n896), .B2(new_n507), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(G1339gat));
  NAND4_X1  g710(.A1(new_n685), .A2(new_n688), .A3(new_n726), .A4(new_n851), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n699), .A2(new_n700), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n711), .A2(new_n712), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n718), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n710), .A2(new_n713), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n708), .B2(new_n701), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n722), .B1(new_n918), .B2(new_n719), .ZN(new_n919));
  INV_X1    g718(.A(new_n723), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n754), .B(new_n916), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n739), .A2(new_n922), .A3(new_n740), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT54), .B1(new_n751), .B2(new_n743), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n735), .A2(new_n743), .A3(new_n738), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n748), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT55), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n751), .A2(new_n743), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n741), .A2(KEYINPUT54), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n930), .A2(KEYINPUT55), .A3(new_n748), .A4(new_n923), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n931), .A3(new_n750), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n921), .B1(new_n932), .B2(new_n726), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n793), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n721), .A2(new_n723), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n630), .A2(new_n935), .A3(new_n916), .ZN(new_n936));
  INV_X1    g735(.A(new_n932), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n913), .B1(new_n939), .B2(new_n684), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(new_n507), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n941), .A2(new_n497), .A3(new_n760), .A4(new_n775), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n259), .A3(new_n726), .ZN(new_n943));
  AOI22_X1  g742(.A1(new_n933), .A2(new_n793), .B1(new_n936), .B2(new_n937), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n912), .B1(new_n944), .B2(new_n686), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n497), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n442), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(new_n760), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n850), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n943), .B1(new_n950), .B2(new_n259), .ZN(G1340gat));
  NOR3_X1   g750(.A1(new_n942), .A2(new_n257), .A3(new_n851), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n754), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n257), .ZN(G1341gat));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n262), .A3(new_n686), .ZN(new_n955));
  OAI21_X1  g754(.A(G127gat), .B1(new_n942), .B2(new_n684), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1342gat));
  NAND2_X1  g756(.A1(new_n760), .A2(new_n630), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n263), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT56), .ZN(new_n961));
  OAI21_X1  g760(.A(G134gat), .B1(new_n942), .B2(new_n793), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(KEYINPUT56), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(G1343gat));
  NOR3_X1   g763(.A1(new_n814), .A2(new_n757), .A3(new_n468), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT57), .B1(new_n940), .B2(new_n500), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT57), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n945), .A2(new_n967), .A3(new_n507), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G141gat), .B1(new_n970), .B2(new_n726), .ZN(new_n971));
  NAND2_X1  g770(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n947), .A2(new_n507), .A3(new_n773), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n973), .A2(new_n468), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n850), .A2(new_n333), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT118), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n971), .A2(new_n972), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g777(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n978), .B(new_n979), .ZN(G1344gat));
  NAND3_X1  g779(.A1(new_n974), .A2(new_n342), .A3(new_n754), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n969), .A3(new_n754), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n342), .A2(KEYINPUT59), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT59), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n985), .B1(new_n982), .B2(G148gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n984), .B2(new_n986), .ZN(G1345gat));
  INV_X1    g786(.A(G155gat), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n970), .A2(new_n988), .A3(new_n684), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n468), .A3(new_n684), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n990), .A2(KEYINPUT120), .ZN(new_n991));
  AOI21_X1  g790(.A(G155gat), .B1(new_n990), .B2(KEYINPUT120), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1346gat));
  OAI21_X1  g792(.A(G162gat), .B1(new_n970), .B2(new_n793), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n959), .A2(new_n618), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n994), .B1(new_n973), .B2(new_n995), .ZN(G1347gat));
  NAND2_X1  g795(.A1(new_n757), .A2(new_n468), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n775), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(new_n941), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n1001), .A2(new_n233), .A3(new_n726), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT121), .ZN(new_n1003));
  INV_X1    g802(.A(new_n442), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n1004), .B2(new_n760), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n442), .A2(KEYINPUT121), .A3(new_n468), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n1005), .A2(new_n757), .A3(new_n945), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT122), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1009), .A2(new_n850), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g810(.A(new_n1002), .B1(new_n1011), .B2(new_n233), .ZN(G1348gat));
  NAND4_X1  g811(.A1(new_n1009), .A2(new_n234), .A3(new_n754), .A4(new_n1010), .ZN(new_n1013));
  OAI21_X1  g812(.A(G176gat), .B1(new_n1001), .B2(new_n851), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1349gat));
  OAI21_X1  g814(.A(G183gat), .B1(new_n1001), .B2(new_n684), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n686), .A2(new_n244), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1016), .B1(new_n1007), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g818(.A1(new_n1009), .A2(new_n247), .A3(new_n630), .A4(new_n1010), .ZN(new_n1020));
  OAI21_X1  g819(.A(G190gat), .B1(new_n1001), .B2(new_n793), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n1021), .A2(KEYINPUT61), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n1021), .A2(KEYINPUT61), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G1351gat));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n966), .A2(new_n968), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n998), .B1(new_n812), .B2(new_n813), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT124), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n773), .A2(KEYINPUT124), .A3(new_n998), .ZN(new_n1030));
  AOI21_X1  g829(.A(new_n1026), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g830(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1025), .B1(new_n1032), .B2(new_n726), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1031), .A2(KEYINPUT125), .A3(new_n850), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n1033), .A2(G197gat), .A3(new_n1034), .ZN(new_n1035));
  NOR3_X1   g834(.A1(new_n1027), .A2(new_n500), .A3(new_n940), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n1036), .A2(new_n372), .A3(new_n850), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1035), .A2(new_n1037), .ZN(G1352gat));
  NAND3_X1  g837(.A1(new_n1036), .A2(new_n373), .A3(new_n754), .ZN(new_n1039));
  XOR2_X1   g838(.A(new_n1039), .B(KEYINPUT62), .Z(new_n1040));
  OAI21_X1  g839(.A(G204gat), .B1(new_n1032), .B2(new_n851), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1040), .A2(new_n1041), .ZN(G1353gat));
  INV_X1    g841(.A(KEYINPUT127), .ZN(new_n1043));
  AOI21_X1  g842(.A(new_n391), .B1(new_n1031), .B2(new_n686), .ZN(new_n1044));
  OAI21_X1  g843(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT63), .ZN(new_n1045));
  AOI21_X1  g844(.A(KEYINPUT124), .B1(new_n773), .B2(new_n998), .ZN(new_n1046));
  AOI211_X1 g845(.A(new_n1028), .B(new_n997), .C1(new_n771), .C2(new_n772), .ZN(new_n1047));
  OAI211_X1 g846(.A(new_n969), .B(new_n686), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g847(.A1(new_n1048), .A2(G211gat), .ZN(new_n1049));
  INV_X1    g848(.A(KEYINPUT63), .ZN(new_n1050));
  NAND3_X1  g849(.A1(new_n1049), .A2(KEYINPUT127), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g850(.A1(new_n1048), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1052));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1053));
  NAND2_X1  g852(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g853(.A1(new_n1048), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1055));
  NAND4_X1  g854(.A1(new_n1045), .A2(new_n1051), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g855(.A1(new_n1036), .A2(new_n391), .A3(new_n686), .ZN(new_n1057));
  NAND2_X1  g856(.A1(new_n1056), .A2(new_n1057), .ZN(G1354gat));
  OAI21_X1  g857(.A(G218gat), .B1(new_n1032), .B2(new_n793), .ZN(new_n1059));
  NAND3_X1  g858(.A1(new_n1036), .A2(new_n392), .A3(new_n630), .ZN(new_n1060));
  NAND2_X1  g859(.A1(new_n1059), .A2(new_n1060), .ZN(G1355gat));
endmodule


