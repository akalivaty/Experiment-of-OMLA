

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U552 ( .A(n527), .B(KEYINPUT65), .ZN(n891) );
  AND2_X1 U553 ( .A1(n778), .A2(n777), .ZN(n519) );
  XOR2_X1 U554 ( .A(KEYINPUT94), .B(n783), .Z(n520) );
  XNOR2_X1 U555 ( .A(KEYINPUT95), .B(n782), .ZN(n521) );
  AND2_X1 U556 ( .A1(n825), .A2(n816), .ZN(n522) );
  AND2_X1 U557 ( .A1(n522), .A2(n817), .ZN(n523) );
  XNOR2_X1 U558 ( .A(KEYINPUT29), .B(KEYINPUT97), .ZN(n524) );
  OR2_X1 U559 ( .A1(n731), .A2(G301), .ZN(n525) );
  INV_X1 U560 ( .A(KEYINPUT96), .ZN(n705) );
  AND2_X1 U561 ( .A1(n730), .A2(n525), .ZN(n740) );
  INV_X1 U562 ( .A(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U563 ( .A1(G8), .A2(n732), .ZN(n781) );
  INV_X1 U564 ( .A(G2104), .ZN(n530) );
  NAND2_X1 U565 ( .A1(G160), .A2(G40), .ZN(n783) );
  NOR2_X1 U566 ( .A1(G651), .A2(n633), .ZN(n655) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n657) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n526), .Z(n887) );
  NAND2_X1 U570 ( .A1(G137), .A2(n887), .ZN(n529) );
  NAND2_X1 U571 ( .A1(n530), .A2(G2105), .ZN(n527) );
  NAND2_X1 U572 ( .A1(G125), .A2(n891), .ZN(n528) );
  NAND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U574 ( .A1(G2105), .A2(n530), .ZN(n549) );
  NAND2_X1 U575 ( .A1(G101), .A2(n549), .ZN(n531) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(n531), .Z(n533) );
  AND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U578 ( .A1(n890), .A2(G113), .ZN(n532) );
  NAND2_X1 U579 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U580 ( .A1(n535), .A2(n534), .ZN(G160) );
  XOR2_X1 U581 ( .A(KEYINPUT104), .B(G2443), .Z(n537) );
  XNOR2_X1 U582 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U583 ( .A(n537), .B(n536), .ZN(n547) );
  XOR2_X1 U584 ( .A(G2427), .B(G2435), .Z(n539) );
  XNOR2_X1 U585 ( .A(G2430), .B(G2438), .ZN(n538) );
  XNOR2_X1 U586 ( .A(n539), .B(n538), .ZN(n543) );
  XOR2_X1 U587 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n541) );
  XNOR2_X1 U588 ( .A(G2446), .B(G2454), .ZN(n540) );
  XNOR2_X1 U589 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U590 ( .A(n543), .B(n542), .Z(n545) );
  XNOR2_X1 U591 ( .A(G2451), .B(KEYINPUT105), .ZN(n544) );
  XNOR2_X1 U592 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U593 ( .A(n547), .B(n546), .ZN(n548) );
  AND2_X1 U594 ( .A1(n548), .A2(G14), .ZN(G401) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U596 ( .A(n549), .Z(n886) );
  NAND2_X1 U597 ( .A1(n886), .A2(G99), .ZN(n550) );
  XOR2_X1 U598 ( .A(KEYINPUT75), .B(n550), .Z(n552) );
  NAND2_X1 U599 ( .A1(n890), .A2(G111), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U601 ( .A(KEYINPUT76), .B(n553), .ZN(n556) );
  NAND2_X1 U602 ( .A1(n891), .A2(G123), .ZN(n554) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(n554), .Z(n555) );
  NOR2_X1 U604 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U605 ( .A1(n887), .A2(G135), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n558), .A2(n557), .ZN(n928) );
  XNOR2_X1 U607 ( .A(G2096), .B(n928), .ZN(n559) );
  OR2_X1 U608 ( .A1(G2100), .A2(n559), .ZN(G156) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G651), .ZN(n564) );
  NOR2_X1 U611 ( .A1(G543), .A2(n564), .ZN(n560) );
  XOR2_X1 U612 ( .A(KEYINPUT1), .B(n560), .Z(n660) );
  NAND2_X1 U613 ( .A1(G64), .A2(n660), .ZN(n562) );
  XOR2_X1 U614 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U615 ( .A1(G52), .A2(n655), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n570) );
  NAND2_X1 U617 ( .A1(n657), .A2(G90), .ZN(n563) );
  XNOR2_X1 U618 ( .A(KEYINPUT67), .B(n563), .ZN(n567) );
  NOR2_X1 U619 ( .A1(n633), .A2(n564), .ZN(n661) );
  NAND2_X1 U620 ( .A1(n661), .A2(G77), .ZN(n565) );
  XOR2_X1 U621 ( .A(KEYINPUT68), .B(n565), .Z(n566) );
  NOR2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U623 ( .A(n568), .B(KEYINPUT9), .ZN(n569) );
  NOR2_X1 U624 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n571), .Z(G171) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  NAND2_X1 U627 ( .A1(n657), .A2(G89), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U629 ( .A1(G76), .A2(n661), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U631 ( .A(n575), .B(KEYINPUT5), .ZN(n581) );
  NAND2_X1 U632 ( .A1(n660), .A2(G63), .ZN(n576) );
  XNOR2_X1 U633 ( .A(n576), .B(KEYINPUT74), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G51), .A2(n655), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U636 ( .A(KEYINPUT6), .B(n579), .Z(n580) );
  NAND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U638 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U640 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n584) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U642 ( .A(n584), .B(n583), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n835) );
  NAND2_X1 U644 ( .A1(n835), .A2(G567), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U646 ( .A1(n660), .A2(G56), .ZN(n586) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n586), .Z(n592) );
  NAND2_X1 U648 ( .A1(n657), .A2(G81), .ZN(n587) );
  XNOR2_X1 U649 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G68), .A2(n661), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U652 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U654 ( .A(n593), .B(KEYINPUT72), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G43), .A2(n655), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n595), .A2(n594), .ZN(n985) );
  INV_X1 U657 ( .A(G860), .ZN(n615) );
  OR2_X1 U658 ( .A1(n985), .A2(n615), .ZN(G153) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U660 ( .A1(G66), .A2(n660), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G92), .A2(n657), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U663 ( .A1(G54), .A2(n655), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G79), .A2(n661), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U666 ( .A(KEYINPUT73), .B(n600), .Z(n601) );
  NOR2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U668 ( .A(KEYINPUT15), .B(n603), .ZN(n976) );
  INV_X1 U669 ( .A(G868), .ZN(n675) );
  NAND2_X1 U670 ( .A1(n976), .A2(n675), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G91), .A2(n657), .ZN(n607) );
  NAND2_X1 U673 ( .A1(G78), .A2(n661), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U675 ( .A1(G65), .A2(n660), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G53), .A2(n655), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U679 ( .A(KEYINPUT70), .B(n612), .Z(G299) );
  NOR2_X1 U680 ( .A1(G299), .A2(G868), .ZN(n614) );
  NOR2_X1 U681 ( .A1(G286), .A2(n675), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n614), .A2(n613), .ZN(G297) );
  NAND2_X1 U683 ( .A1(n615), .A2(G559), .ZN(n616) );
  INV_X1 U684 ( .A(n976), .ZN(n627) );
  NAND2_X1 U685 ( .A1(n616), .A2(n627), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n617), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n985), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n627), .A2(G868), .ZN(n618) );
  NOR2_X1 U689 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G93), .A2(n657), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G80), .A2(n661), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G67), .A2(n660), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G55), .A2(n655), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n674) );
  NAND2_X1 U698 ( .A1(G559), .A2(n627), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(n985), .ZN(n672) );
  XOR2_X1 U700 ( .A(n672), .B(KEYINPUT77), .Z(n629) );
  NOR2_X1 U701 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U702 ( .A(KEYINPUT78), .B(n630), .Z(n631) );
  XNOR2_X1 U703 ( .A(n674), .B(n631), .ZN(G145) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(KEYINPUT80), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n633), .A2(G87), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U708 ( .A1(n660), .A2(n636), .ZN(n639) );
  NAND2_X1 U709 ( .A1(G49), .A2(n655), .ZN(n637) );
  XOR2_X1 U710 ( .A(KEYINPUT79), .B(n637), .Z(n638) );
  NAND2_X1 U711 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G60), .A2(n660), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G47), .A2(n655), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT66), .B(n642), .Z(n646) );
  NAND2_X1 U716 ( .A1(G85), .A2(n657), .ZN(n644) );
  NAND2_X1 U717 ( .A1(G72), .A2(n661), .ZN(n643) );
  AND2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G73), .A2(n661), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT2), .ZN(n654) );
  NAND2_X1 U722 ( .A1(G61), .A2(n660), .ZN(n649) );
  NAND2_X1 U723 ( .A1(G48), .A2(n655), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G86), .A2(n657), .ZN(n650) );
  XNOR2_X1 U726 ( .A(KEYINPUT81), .B(n650), .ZN(n651) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U729 ( .A1(n655), .A2(G50), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT82), .ZN(n659) );
  NAND2_X1 U731 ( .A1(G88), .A2(n657), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n665) );
  NAND2_X1 U733 ( .A1(G62), .A2(n660), .ZN(n663) );
  NAND2_X1 U734 ( .A1(G75), .A2(n661), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U736 ( .A1(n665), .A2(n664), .ZN(G166) );
  XOR2_X1 U737 ( .A(G290), .B(G305), .Z(n666) );
  XNOR2_X1 U738 ( .A(G288), .B(n666), .ZN(n669) );
  XOR2_X1 U739 ( .A(n674), .B(KEYINPUT19), .Z(n667) );
  XNOR2_X1 U740 ( .A(n667), .B(KEYINPUT83), .ZN(n668) );
  XOR2_X1 U741 ( .A(n669), .B(n668), .Z(n671) );
  XNOR2_X1 U742 ( .A(G166), .B(G299), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n905) );
  XNOR2_X1 U744 ( .A(n672), .B(n905), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n673), .A2(G868), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n681), .A2(G2072), .ZN(n682) );
  XNOR2_X1 U753 ( .A(KEYINPUT84), .B(n682), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U755 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n684) );
  NAND2_X1 U756 ( .A1(G132), .A2(G82), .ZN(n683) );
  XNOR2_X1 U757 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U758 ( .A1(n685), .A2(G218), .ZN(n686) );
  NAND2_X1 U759 ( .A1(G96), .A2(n686), .ZN(n840) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n840), .ZN(n690) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n687) );
  NOR2_X1 U762 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U763 ( .A1(G108), .A2(n688), .ZN(n841) );
  NAND2_X1 U764 ( .A1(G567), .A2(n841), .ZN(n689) );
  NAND2_X1 U765 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U766 ( .A(KEYINPUT86), .B(n691), .Z(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n693) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U769 ( .A1(n693), .A2(n692), .ZN(n839) );
  NAND2_X1 U770 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U771 ( .A1(G102), .A2(n886), .ZN(n695) );
  NAND2_X1 U772 ( .A1(G138), .A2(n887), .ZN(n694) );
  NAND2_X1 U773 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U774 ( .A1(G114), .A2(n890), .ZN(n697) );
  NAND2_X1 U775 ( .A1(G126), .A2(n891), .ZN(n696) );
  NAND2_X1 U776 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U777 ( .A1(n699), .A2(n698), .ZN(G164) );
  INV_X1 U778 ( .A(G166), .ZN(G303) );
  XOR2_X1 U779 ( .A(G1981), .B(G305), .Z(n968) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n784) );
  AND2_X1 U781 ( .A1(n784), .A2(n520), .ZN(n727) );
  INV_X1 U782 ( .A(n727), .ZN(n732) );
  AND2_X1 U783 ( .A1(G1341), .A2(n732), .ZN(n700) );
  NOR2_X1 U784 ( .A1(n985), .A2(n700), .ZN(n704) );
  NAND2_X1 U785 ( .A1(n727), .A2(G1996), .ZN(n702) );
  XOR2_X1 U786 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n701) );
  XOR2_X1 U787 ( .A(n702), .B(n701), .Z(n703) );
  NAND2_X1 U788 ( .A1(n704), .A2(n703), .ZN(n716) );
  NOR2_X1 U789 ( .A1(n716), .A2(n976), .ZN(n706) );
  XNOR2_X1 U790 ( .A(n706), .B(n705), .ZN(n714) );
  NOR2_X1 U791 ( .A1(n727), .A2(G1348), .ZN(n708) );
  NOR2_X1 U792 ( .A1(G2067), .A2(n732), .ZN(n707) );
  NOR2_X1 U793 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n727), .A2(G2072), .ZN(n709) );
  XNOR2_X1 U795 ( .A(n709), .B(KEYINPUT27), .ZN(n711) );
  INV_X1 U796 ( .A(G1956), .ZN(n992) );
  NOR2_X1 U797 ( .A1(n992), .A2(n727), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n720) );
  INV_X1 U799 ( .A(G299), .ZN(n719) );
  NAND2_X1 U800 ( .A1(n720), .A2(n719), .ZN(n715) );
  AND2_X1 U801 ( .A1(n712), .A2(n715), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n725) );
  INV_X1 U803 ( .A(n715), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n716), .A2(n976), .ZN(n717) );
  OR2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n723) );
  NOR2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U807 ( .A(n721), .B(KEYINPUT28), .Z(n722) );
  AND2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U810 ( .A(n726), .B(n524), .ZN(n730) );
  XOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NOR2_X1 U812 ( .A1(n948), .A2(n732), .ZN(n729) );
  NOR2_X1 U813 ( .A1(n727), .A2(G1961), .ZN(n728) );
  NOR2_X1 U814 ( .A1(n729), .A2(n728), .ZN(n731) );
  AND2_X1 U815 ( .A1(G301), .A2(n731), .ZN(n737) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n781), .ZN(n757) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n732), .ZN(n753) );
  NOR2_X1 U818 ( .A1(n757), .A2(n753), .ZN(n733) );
  NAND2_X1 U819 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G168), .A2(n735), .ZN(n736) );
  NOR2_X1 U822 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U823 ( .A(n738), .B(KEYINPUT31), .ZN(n739) );
  NOR2_X1 U824 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U825 ( .A(n742), .B(n741), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n755), .A2(G286), .ZN(n750) );
  INV_X1 U827 ( .A(G8), .ZN(n748) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n781), .ZN(n744) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n732), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U831 ( .A(KEYINPUT99), .B(n745), .Z(n746) );
  NAND2_X1 U832 ( .A1(n746), .A2(G303), .ZN(n747) );
  OR2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n749) );
  AND2_X1 U834 ( .A1(n750), .A2(n749), .ZN(n752) );
  XOR2_X1 U835 ( .A(KEYINPUT100), .B(KEYINPUT32), .Z(n751) );
  XNOR2_X1 U836 ( .A(n752), .B(n751), .ZN(n759) );
  NAND2_X1 U837 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U839 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U840 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U841 ( .A(n760), .B(KEYINPUT101), .ZN(n775) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NOR2_X1 U844 ( .A1(n761), .A2(n973), .ZN(n763) );
  INV_X1 U845 ( .A(KEYINPUT33), .ZN(n762) );
  AND2_X1 U846 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U847 ( .A1(n775), .A2(n764), .ZN(n768) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U849 ( .A(n974), .ZN(n765) );
  NOR2_X1 U850 ( .A1(n765), .A2(n781), .ZN(n766) );
  OR2_X1 U851 ( .A1(KEYINPUT33), .A2(n766), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U853 ( .A1(n973), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U854 ( .A1(n769), .A2(n781), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n968), .A2(n772), .ZN(n778) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n776), .A2(n781), .ZN(n777) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U862 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  NOR2_X1 U863 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U864 ( .A1(n519), .A2(n521), .ZN(n818) );
  NOR2_X1 U865 ( .A1(n784), .A2(n783), .ZN(n829) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NAND2_X1 U867 ( .A1(n887), .A2(G140), .ZN(n785) );
  XOR2_X1 U868 ( .A(KEYINPUT87), .B(n785), .Z(n787) );
  NAND2_X1 U869 ( .A1(n886), .A2(G104), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n788), .ZN(n794) );
  NAND2_X1 U872 ( .A1(G116), .A2(n890), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G128), .A2(n891), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U875 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  XNOR2_X1 U876 ( .A(KEYINPUT88), .B(n792), .ZN(n793) );
  NOR2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U878 ( .A(n795), .B(KEYINPUT36), .Z(n796) );
  XNOR2_X1 U879 ( .A(KEYINPUT89), .B(n796), .ZN(n902) );
  NOR2_X1 U880 ( .A1(n827), .A2(n902), .ZN(n939) );
  NAND2_X1 U881 ( .A1(n829), .A2(n939), .ZN(n825) );
  XNOR2_X1 U882 ( .A(n829), .B(KEYINPUT92), .ZN(n814) );
  NAND2_X1 U883 ( .A1(G117), .A2(n890), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G129), .A2(n891), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n886), .A2(G105), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n887), .A2(G141), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n881) );
  NAND2_X1 U891 ( .A1(G1996), .A2(n881), .ZN(n804) );
  XOR2_X1 U892 ( .A(KEYINPUT91), .B(n804), .Z(n813) );
  NAND2_X1 U893 ( .A1(G95), .A2(n886), .ZN(n806) );
  NAND2_X1 U894 ( .A1(G107), .A2(n890), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n891), .A2(G119), .ZN(n807) );
  XOR2_X1 U897 ( .A(KEYINPUT90), .B(n807), .Z(n808) );
  NOR2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n887), .A2(G131), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n811), .A2(n810), .ZN(n897) );
  NAND2_X1 U901 ( .A1(G1991), .A2(n897), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n927) );
  NAND2_X1 U903 ( .A1(n814), .A2(n927), .ZN(n815) );
  XNOR2_X1 U904 ( .A(n815), .B(KEYINPUT93), .ZN(n822) );
  INV_X1 U905 ( .A(n822), .ZN(n816) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U907 ( .A1(n982), .A2(n829), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n523), .ZN(n832) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n881), .ZN(n931) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n897), .ZN(n923) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n819) );
  XNOR2_X1 U912 ( .A(KEYINPUT102), .B(n819), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n923), .A2(n820), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U915 ( .A1(n931), .A2(n823), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n824), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n827), .A2(n902), .ZN(n936) );
  NAND2_X1 U919 ( .A1(n828), .A2(n936), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U922 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n833) );
  XNOR2_X1 U923 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n836) );
  XOR2_X1 U926 ( .A(KEYINPUT108), .B(n836), .Z(n837) );
  NAND2_X1 U927 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2090), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2084), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n844), .B(G2100), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2078), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2678), .B(KEYINPUT109), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n850), .B(n849), .Z(G227) );
  XOR2_X1 U948 ( .A(KEYINPUT111), .B(G1961), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1971), .B(G1956), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G1966), .B(G1976), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1981), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT110), .B(G2474), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U960 ( .A1(n891), .A2(G124), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G136), .A2(n887), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(KEYINPUT112), .B(n865), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G100), .A2(n886), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G112), .A2(n890), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G118), .A2(n890), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G130), .A2(n891), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G106), .A2(n886), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G142), .A2(n887), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(n928), .ZN(n885) );
  XOR2_X1 U978 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n879) );
  XNOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U982 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n899) );
  NAND2_X1 U985 ( .A1(G103), .A2(n886), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G139), .A2(n887), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U988 ( .A1(G115), .A2(n890), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n916) );
  XNOR2_X1 U993 ( .A(n897), .B(n916), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(G162), .B(n900), .Z(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U998 ( .A(KEYINPUT115), .B(n976), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n904), .B(n985), .ZN(n906) );
  XOR2_X1 U1000 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1001 ( .A(G286), .B(G171), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1005 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  NAND2_X1 U1006 ( .A1(n911), .A2(G319), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(KEYINPUT116), .B(n913), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1013 ( .A(G2072), .B(n916), .Z(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT118), .B(n917), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(G2078), .B(G164), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(KEYINPUT119), .B(n918), .ZN(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT50), .B(n921), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n932), .Z(n933) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(n933), .ZN(n934) );
  NOR2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  XOR2_X1 U1032 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n963) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n963), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n942), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G35), .ZN(n957) );
  XNOR2_X1 U1036 ( .A(G1996), .B(G32), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT121), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(n951), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G25), .B(G1991), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n955), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(n958), .Z(n961) );
  XOR2_X1 U1051 ( .A(KEYINPUT54), .B(G34), .Z(n959) );
  XNOR2_X1 U1052 ( .A(G2084), .B(n959), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1055 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n966), .ZN(n1020) );
  INV_X1 U1058 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1059 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n967) );
  XNOR2_X1 U1060 ( .A(n1016), .B(n967), .ZN(n991) );
  XNOR2_X1 U1061 ( .A(G168), .B(G1966), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n970), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1064 ( .A(G171), .B(G1961), .ZN(n984) );
  XNOR2_X1 U1065 ( .A(G303), .B(G1971), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT125), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(G1956), .B(G299), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1348), .B(n976), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n985), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n1018) );
  XNOR2_X1 U1079 ( .A(G20), .B(n992), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G1981), .B(G6), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G19), .B(G1341), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1084 ( .A(KEYINPUT59), .B(G1348), .Z(n997) );
  XNOR2_X1 U1085 ( .A(G4), .B(n997), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT60), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1088 ( .A(G1961), .B(G5), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1012) );
  XNOR2_X1 U1090 ( .A(G1966), .B(KEYINPUT126), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1003), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G1976), .B(G23), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT127), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

