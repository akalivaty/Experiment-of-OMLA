//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI211_X1 g009(.A(KEYINPUT1), .B(G127gat), .C1(new_n205), .C2(new_n207), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n202), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G141gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G155gat), .B(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT2), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231));
  OAI21_X1  g030(.A(G127gat), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n208), .A2(new_n209), .A3(new_n203), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(G134gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n212), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT4), .ZN(new_n236));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n229), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT75), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n219), .A2(new_n229), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n241), .A2(new_n244), .B1(new_n212), .B2(new_n234), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n236), .A2(new_n239), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n212), .A2(new_n234), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n235), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n252), .B2(new_n238), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n256), .B1(new_n246), .B2(new_n245), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G1gat), .B(G29gat), .Z(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n236), .A2(new_n247), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n238), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n270), .B(KEYINPUT39), .C1(new_n238), .C2(new_n252), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT39), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n272), .A3(new_n238), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT80), .A3(new_n265), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT80), .B1(new_n273), .B2(new_n265), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT40), .B(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n268), .B1(new_n277), .B2(KEYINPUT81), .ZN(new_n278));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(G169gat), .ZN(new_n288));
  INV_X1    g087(.A(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n279), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n290), .A2(new_n291), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n307));
  OR2_X1    g106(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n309));
  AOI21_X1  g108(.A(G190gat), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n310), .B2(KEYINPUT65), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT26), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n293), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n279), .C1(new_n315), .C2(new_n312), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n307), .ZN(new_n318));
  INV_X1    g117(.A(new_n309), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n284), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n311), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G211gat), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G211gat), .A2(G218gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n338));
  AND2_X1   g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n343), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT69), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n337), .B(new_n338), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n336), .A2(new_n345), .A3(new_n346), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(KEYINPUT69), .A3(new_n346), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n337), .A4(new_n338), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n349), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n329), .A2(new_n331), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n349), .A2(new_n350), .A3(new_n355), .ZN(new_n358));
  INV_X1    g157(.A(new_n331), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n330), .B1(new_n325), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(KEYINPUT74), .B(G36gat), .Z(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT73), .B(G8gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n357), .A2(new_n362), .A3(new_n368), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n363), .A2(new_n373), .A3(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n276), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n274), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT40), .A4(new_n271), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT40), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n278), .A2(new_n376), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n248), .A2(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT6), .B1(new_n385), .B2(new_n265), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n267), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n260), .A2(KEYINPUT6), .A3(new_n266), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n329), .A2(new_n331), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n358), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n359), .A2(new_n361), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n392), .B(KEYINPUT37), .C1(new_n393), .C2(new_n358), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT37), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT82), .B1(new_n363), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n397), .B(KEYINPUT37), .C1(new_n357), .C2(new_n362), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n394), .B(new_n368), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT38), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n399), .A2(new_n400), .A3(new_n370), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n396), .A2(new_n398), .B1(new_n395), .B2(new_n363), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n402), .A2(new_n400), .A3(new_n369), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n390), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n326), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n241), .B2(new_n244), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n356), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n358), .B2(new_n360), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n408), .B(new_n410), .C1(new_n411), .C2(new_n230), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n335), .B(new_n334), .C1(new_n341), .C2(new_n343), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n350), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n240), .A3(new_n326), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n246), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT77), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n418), .A3(new_n246), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n417), .B(new_n419), .C1(new_n358), .C2(new_n406), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n409), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  INV_X1    g222(.A(G22gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(G78gat), .B(G106gat), .Z(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT31), .ZN(new_n428));
  INV_X1    g227(.A(G50gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n412), .B(new_n421), .C1(new_n423), .C2(new_n424), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n426), .A2(KEYINPUT79), .A3(new_n431), .A4(new_n430), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n422), .A2(new_n424), .ZN(new_n436));
  INV_X1    g235(.A(new_n430), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n412), .A2(G22gat), .A3(new_n421), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n384), .A2(new_n404), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n311), .A2(new_n317), .A3(new_n323), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n295), .B1(new_n300), .B2(new_n302), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n304), .A2(new_n443), .B1(new_n294), .B2(new_n295), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n250), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n306), .A2(new_n234), .A3(new_n324), .A4(new_n212), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G227gat), .ZN(new_n448));
  INV_X1    g247(.A(G233gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT67), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT67), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n452), .B(new_n453), .C1(new_n445), .C2(new_n446), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT32), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g256(.A(G15gat), .B(G43gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  OAI221_X1 g261(.A(KEYINPUT32), .B1(new_n456), .B2(new_n462), .C1(new_n451), .C2(new_n454), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n453), .A3(new_n446), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT34), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g267(.A(new_n466), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n461), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n461), .B2(new_n463), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(KEYINPUT36), .A3(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n461), .A2(new_n469), .A3(new_n463), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n440), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n389), .A2(new_n375), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n441), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n387), .A2(new_n388), .B1(new_n374), .B2(new_n372), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n475), .A2(new_n472), .A3(KEYINPUT68), .ZN(new_n486));
  INV_X1    g285(.A(new_n473), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n440), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n440), .A2(new_n490), .A3(new_n476), .A4(new_n485), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G57gat), .B(G64gat), .Z(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(KEYINPUT9), .ZN(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G78gat), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(KEYINPUT88), .A2(G64gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT88), .A2(G64gat), .ZN(new_n499));
  OAI21_X1  g298(.A(G57gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n502), .B(KEYINPUT90), .Z(new_n503));
  INV_X1    g302(.A(G64gat), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n500), .B(KEYINPUT89), .C1(G57gat), .C2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(new_n503), .A3(new_n505), .A4(new_n496), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G15gat), .B(G22gat), .Z(new_n513));
  INV_X1    g312(.A(G1gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n518), .A3(KEYINPUT85), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(G8gat), .C1(KEYINPUT85), .C2(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT86), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n522), .A2(new_n523), .A3(G8gat), .A4(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G8gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n518), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT87), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n525), .B(new_n528), .C1(new_n508), .C2(new_n507), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(G183gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(G183gat), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n533), .ZN(new_n537));
  XNOR2_X1  g336(.A(G127gat), .B(G155gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(new_n332), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n535), .B2(new_n537), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n512), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n535), .A2(new_n537), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n511), .A3(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550));
  INV_X1    g349(.A(G43gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(G50gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n552), .B2(KEYINPUT84), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT14), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n555), .A2(G29gat), .A3(G36gat), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n557), .A2(new_n556), .A3(new_n554), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n558), .B(new_n559), .C1(new_n561), .C2(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT17), .ZN(new_n564));
  XOR2_X1   g363(.A(G99gat), .B(G106gat), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT92), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT91), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT7), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n567), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n569), .A2(new_n575), .A3(new_n565), .A4(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT93), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n563), .A2(new_n579), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n585), .A3(new_n580), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n582), .A2(new_n590), .A3(new_n584), .A4(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n595), .A3(new_n591), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n493), .A2(new_n549), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n507), .A2(new_n579), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n574), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n565), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n574), .A2(new_n603), .A3(new_n566), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(new_n506), .A3(new_n497), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT95), .B(KEYINPUT10), .Z(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n602), .B2(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n579), .A2(KEYINPUT10), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n507), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n609), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n608), .A2(KEYINPUT96), .A3(new_n609), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n289), .ZN(new_n621));
  INV_X1    g420(.A(G204gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n617), .A2(new_n623), .A3(new_n618), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n525), .A2(new_n528), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n563), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n563), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT17), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n563), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n633), .A2(new_n525), .A3(new_n528), .A4(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n631), .B(KEYINPUT13), .Z(new_n640));
  NOR2_X1   g439(.A1(new_n629), .A2(new_n563), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n632), .B1(new_n525), .B2(new_n528), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n630), .A2(new_n636), .A3(KEYINPUT18), .A4(new_n631), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(G169gat), .B(G197gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n639), .A2(new_n643), .A3(new_n644), .A4(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n601), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n389), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n514), .ZN(G1324gat));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT97), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n658), .A2(new_n375), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n665), .B2(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI211_X1 g468(.A(KEYINPUT97), .B(new_n661), .C1(new_n663), .C2(new_n664), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n669), .A2(new_n670), .B1(new_n526), .B2(new_n663), .ZN(G1325gat));
  INV_X1    g470(.A(new_n658), .ZN(new_n672));
  AOI21_X1  g471(.A(G15gat), .B1(new_n672), .B2(new_n476), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n479), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n474), .A2(KEYINPUT99), .A3(new_n478), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT100), .Z(new_n679));
  AOI21_X1  g478(.A(new_n673), .B1(new_n672), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n658), .A2(new_n440), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n493), .A2(new_n599), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n548), .A2(new_n628), .A3(new_n656), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(G29gat), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(KEYINPUT102), .A3(new_n687), .A4(new_n390), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(new_n390), .A3(new_n685), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(G29gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n492), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n489), .A2(KEYINPUT104), .A3(new_n491), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n434), .A2(new_n435), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n698), .A2(KEYINPUT103), .A3(new_n482), .A4(new_n439), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n440), .B2(new_n485), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n675), .A2(new_n441), .A3(new_n702), .A4(new_n676), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n697), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n600), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n493), .B2(new_n599), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n685), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n389), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT105), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n694), .B1(new_n711), .B2(new_n687), .ZN(G1328gat));
  INV_X1    g511(.A(new_n686), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(G36gat), .A3(new_n375), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  OAI21_X1  g514(.A(G36gat), .B1(new_n709), .B2(new_n375), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(new_n476), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n713), .A2(G43gat), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n708), .A2(new_n685), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n677), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n721), .B2(new_n677), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT47), .B(new_n720), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n551), .B1(new_n721), .B2(new_n677), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n719), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(G1330gat));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  OAI21_X1  g530(.A(G50gat), .B1(new_n709), .B2(new_n440), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n686), .A2(new_n429), .A3(new_n481), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(KEYINPUT107), .A3(new_n733), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT107), .B2(new_n732), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(new_n731), .ZN(G1331gat));
  NOR3_X1   g536(.A1(new_n549), .A2(new_n655), .A3(new_n600), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n704), .A2(new_n628), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n390), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n376), .B1(new_n748), .B2(new_n504), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT109), .Z(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n744), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT110), .B1(new_n743), .B2(new_n750), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n504), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n752), .A2(new_n748), .A3(new_n753), .A4(new_n504), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n744), .A2(G71gat), .A3(new_n677), .ZN(new_n759));
  INV_X1    g558(.A(G71gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n743), .B2(new_n718), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT50), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n744), .A2(new_n481), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n548), .A2(new_n655), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n706), .B2(new_n707), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n628), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n772), .A2(new_n571), .A3(new_n389), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n704), .A2(new_n600), .A3(new_n769), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n600), .A4(new_n769), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n627), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n390), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n773), .A2(new_n779), .ZN(G1336gat));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n772), .A2(new_n572), .A3(new_n375), .ZN(new_n782));
  AOI21_X1  g581(.A(G92gat), .B1(new_n778), .B2(new_n376), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n781), .B(new_n786), .C1(new_n782), .C2(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1337gat));
  INV_X1    g587(.A(new_n677), .ZN(new_n789));
  OAI21_X1  g588(.A(G99gat), .B1(new_n772), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n776), .A2(new_n777), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n718), .A2(G99gat), .A3(new_n627), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT112), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n792), .B2(new_n794), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n708), .A2(new_n628), .A3(new_n481), .A4(new_n769), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT113), .B(G106gat), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n771), .A2(new_n799), .A3(new_n628), .A4(new_n481), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n791), .A2(new_n803), .A3(new_n628), .A4(new_n481), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n796), .A2(new_n798), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n804), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n808), .B2(KEYINPUT53), .ZN(new_n809));
  AOI211_X1 g608(.A(KEYINPUT114), .B(new_n802), .C1(new_n807), .C2(new_n804), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n805), .B1(new_n809), .B2(new_n810), .ZN(G1339gat));
  NOR3_X1   g610(.A1(new_n612), .A2(new_n609), .A3(new_n614), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n615), .B1(new_n812), .B2(KEYINPUT116), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n611), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n608), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n614), .ZN(new_n817));
  INV_X1    g616(.A(new_n609), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT116), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT54), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n624), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n818), .B1(new_n816), .B2(new_n817), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n822), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n623), .B(new_n825), .C1(new_n813), .C2(new_n820), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n626), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n826), .A2(new_n830), .A3(new_n831), .A4(new_n655), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n641), .A2(new_n642), .A3(new_n640), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n631), .B1(new_n630), .B2(new_n636), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n650), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n654), .B(new_n835), .C1(new_n625), .C2(new_n626), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n832), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n599), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n826), .A2(new_n830), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n654), .A2(new_n835), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n597), .A2(new_n598), .B1(KEYINPUT118), .B2(new_n843), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n842), .A2(new_n844), .A3(new_n845), .A4(new_n831), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n548), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n627), .A2(new_n548), .A3(new_n656), .A4(new_n599), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(new_n718), .A3(new_n481), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n389), .A2(new_n376), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n656), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n847), .A2(new_n848), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n486), .A2(new_n487), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n481), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n854), .A2(new_n855), .A3(new_n390), .A4(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n390), .B(new_n857), .C1(new_n847), .C2(new_n848), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT120), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n375), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n655), .A2(new_n206), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT121), .Z(new_n863));
  OAI21_X1  g662(.A(new_n853), .B1(new_n861), .B2(new_n863), .ZN(G1340gat));
  OR3_X1    g663(.A1(new_n861), .A2(G120gat), .A3(new_n627), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n852), .B2(new_n627), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  OAI21_X1  g666(.A(new_n203), .B1(new_n861), .B2(new_n549), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n850), .A2(G127gat), .A3(new_n548), .A4(new_n851), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT122), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1342gat));
  NAND2_X1  g673(.A1(new_n600), .A2(new_n202), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n861), .A2(KEYINPUT56), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n852), .B2(new_n599), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT56), .B1(new_n861), .B2(new_n875), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n789), .A2(new_n851), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n837), .A2(new_n599), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n548), .B1(new_n881), .B2(new_n846), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n481), .B1(new_n882), .B2(new_n848), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(new_n481), .C1(new_n847), .C2(new_n848), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n886), .A3(new_n655), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n849), .A2(new_n440), .ZN(new_n889));
  INV_X1    g688(.A(new_n880), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n889), .A2(new_n220), .A3(new_n655), .A4(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n888), .B2(new_n891), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n888), .A2(new_n891), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT123), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT58), .B1(new_n899), .B2(new_n893), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n897), .A2(new_n900), .ZN(G1344gat));
  NAND4_X1  g700(.A1(new_n889), .A2(new_n222), .A3(new_n628), .A4(new_n890), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT124), .Z(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT57), .B(new_n481), .C1(new_n847), .C2(new_n848), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n883), .A2(new_n885), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n628), .A3(new_n890), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n884), .A2(new_n886), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n904), .B1(new_n910), .B2(new_n627), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n222), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n909), .B2(new_n912), .ZN(G1345gat));
  NOR3_X1   g712(.A1(new_n910), .A2(new_n226), .A3(new_n549), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n889), .A2(new_n548), .A3(new_n890), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n226), .B2(new_n915), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n910), .A2(new_n227), .A3(new_n599), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n889), .A2(new_n600), .A3(new_n890), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n227), .B2(new_n918), .ZN(G1347gat));
  NOR3_X1   g718(.A1(new_n849), .A2(new_n856), .A3(new_n481), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n390), .A2(new_n375), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n288), .A3(new_n655), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n850), .A2(new_n921), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n656), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1348gat));
  NOR3_X1   g726(.A1(new_n925), .A2(new_n289), .A3(new_n627), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n628), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n289), .B2(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n925), .B2(new_n549), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n548), .B1(new_n320), .B2(new_n319), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n922), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n931), .B(new_n935), .C1(new_n922), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n923), .A2(new_n284), .A3(new_n600), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n850), .A2(new_n600), .A3(new_n921), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(G190gat), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n939), .B2(G190gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n789), .A2(new_n921), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n889), .A2(new_n946), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n947), .A2(G197gat), .A3(new_n656), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n907), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n656), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1352gat));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n947), .A2(G204gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n628), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n907), .A2(new_n628), .A3(new_n946), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n953), .A2(KEYINPUT125), .A3(new_n959), .A4(new_n628), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n960), .ZN(G1353gat));
  AOI211_X1 g760(.A(new_n549), .B(new_n945), .C1(new_n905), .C2(new_n906), .ZN(new_n962));
  OAI211_X1 g761(.A(KEYINPUT126), .B(KEYINPUT63), .C1(new_n962), .C2(new_n332), .ZN(new_n963));
  INV_X1    g762(.A(new_n947), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n332), .A3(new_n548), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n907), .A2(new_n548), .A3(new_n946), .ZN(new_n966));
  NAND2_X1  g765(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n967));
  OR2_X1    g766(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n966), .A2(G211gat), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n963), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n963), .A2(new_n972), .A3(new_n969), .A4(new_n965), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1354gat));
  NAND3_X1  g773(.A1(new_n964), .A2(new_n333), .A3(new_n600), .ZN(new_n975));
  OAI21_X1  g774(.A(G218gat), .B1(new_n949), .B2(new_n599), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


