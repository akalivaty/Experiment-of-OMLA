//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n189), .A2(new_n190), .B1(G104), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G104), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n192), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n193), .A2(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n190), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n194), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  INV_X1    g021(.A(G116), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT2), .B(G113), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n210), .A2(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n219), .B(G101), .C1(new_n192), .C2(new_n197), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n205), .A2(new_n217), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n191), .A2(G104), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n201), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n204), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n207), .A2(new_n209), .A3(new_n213), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n213), .B1(new_n207), .B2(new_n209), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT5), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G113), .B1(new_n207), .B2(KEYINPUT5), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n230), .A3(new_n216), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n222), .B1(new_n201), .B2(new_n190), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n203), .B1(new_n233), .B2(new_n200), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n219), .A2(new_n234), .B1(new_n215), .B2(new_n216), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n218), .B1(new_n235), .B2(new_n205), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n188), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n205), .A2(new_n217), .A3(new_n220), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT82), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(new_n187), .A3(new_n231), .A4(new_n221), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n237), .A2(new_n240), .A3(new_n241), .A4(KEYINPUT6), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(new_n188), .C1(new_n232), .C2(new_n236), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT83), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G143), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n248), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT0), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n251), .B2(G146), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(KEYINPUT66), .A3(G143), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n252), .A4(new_n248), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n250), .A2(new_n252), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT68), .A2(G128), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT68), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(G143), .B2(new_n249), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n267), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n262), .A2(new_n263), .A3(new_n274), .A4(new_n252), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n266), .A2(KEYINPUT84), .B1(G125), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n266), .A2(KEYINPUT84), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G224), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(G224), .B(new_n280), .C1(new_n277), .C2(new_n278), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n247), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n281), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n240), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n277), .B2(new_n278), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n204), .A2(new_n223), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n230), .A2(new_n216), .A3(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT5), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n216), .B1(new_n294), .B2(new_n228), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n224), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n187), .B(KEYINPUT8), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n283), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n287), .B1(new_n289), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n285), .A2(new_n286), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n286), .ZN(new_n303));
  INV_X1    g117(.A(new_n284), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT83), .A3(new_n245), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n306), .B2(new_n242), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n307), .B2(new_n300), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n280), .A2(G227), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT78), .ZN(new_n313));
  XNOR2_X1  g127(.A(G110), .B(G140), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  AOI21_X1  g132(.A(G131), .B1(new_n317), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n319), .A3(new_n324), .A4(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n318), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G131), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n273), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT70), .B1(new_n273), .B2(new_n275), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n292), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n265), .B1(new_n219), .B2(new_n234), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n334), .A2(new_n336), .B1(new_n337), .B2(new_n205), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n262), .A2(new_n263), .A3(new_n252), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n251), .A2(G146), .ZN(new_n341));
  OAI21_X1  g155(.A(G128), .B1(new_n341), .B2(new_n271), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AND4_X1   g157(.A1(new_n262), .A2(new_n263), .A3(new_n274), .A4(new_n252), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n204), .B(new_n223), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n339), .B1(new_n345), .B2(new_n335), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n340), .B2(new_n342), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n339), .B(new_n335), .C1(new_n348), .C2(new_n292), .ZN(new_n349));
  AND4_X1   g163(.A1(new_n331), .A2(new_n338), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n346), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n331), .B1(new_n352), .B2(new_n338), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n315), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n331), .A3(new_n338), .ZN(new_n355));
  INV_X1    g169(.A(new_n315), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT81), .B1(new_n224), .B2(new_n276), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n292), .A2(new_n358), .A3(new_n275), .A4(new_n273), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n345), .A3(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n360), .A2(KEYINPUT12), .A3(new_n330), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT12), .B1(new_n360), .B2(new_n330), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n355), .B(new_n356), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G469), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n287), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n355), .B1(new_n361), .B2(new_n362), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n315), .ZN(new_n368));
  INV_X1    g182(.A(new_n353), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n356), .A3(new_n355), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(G469), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n365), .A2(new_n287), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n366), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n311), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n280), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n251), .ZN(new_n381));
  NAND2_X1  g195(.A1(G143), .A2(G214), .ZN(new_n382));
  NOR4_X1   g196(.A1(new_n382), .A2(KEYINPUT85), .A3(G237), .A4(G953), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n384));
  AND2_X1   g198(.A1(G143), .A2(G214), .ZN(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n381), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G140), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G125), .ZN(new_n392));
  INV_X1    g206(.A(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n394), .A3(new_n249), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n388), .B2(new_n389), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT75), .A4(KEYINPUT16), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT16), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n392), .B2(KEYINPUT16), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G146), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(KEYINPUT17), .A3(G131), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n249), .B(new_n401), .C1(new_n402), .C2(new_n404), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(G131), .B1(new_n380), .B2(new_n251), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n387), .B2(new_n383), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT86), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n388), .A2(G131), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT17), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n410), .B(new_n415), .C1(new_n387), .C2(new_n383), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n412), .A2(new_n413), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n400), .B1(new_n409), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G113), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n193), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT87), .Z(new_n421));
  OR2_X1    g235(.A1(new_n388), .A2(new_n389), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n388), .A2(new_n389), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n398), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n412), .A2(new_n413), .A3(new_n416), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n395), .B(KEYINPUT19), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n406), .B1(new_n426), .B2(G146), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n420), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n418), .A2(new_n421), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G475), .A2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT20), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n409), .A2(new_n417), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n424), .A3(new_n421), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n429), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n431), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n434), .A2(new_n424), .A3(new_n421), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n418), .A2(new_n420), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n287), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G475), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G952), .ZN(new_n446));
  AOI211_X1 g260(.A(G953), .B(new_n446), .C1(G234), .C2(G237), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n287), .B(new_n280), .C1(G234), .C2(G237), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(G898), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(KEYINPUT68), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT68), .A2(G128), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(G143), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT13), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n256), .A2(G143), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n456), .A2(G134), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n454), .A2(KEYINPUT13), .A3(G134), .A4(new_n458), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT88), .B1(new_n208), .B2(G122), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n463));
  INV_X1    g277(.A(G122), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(G116), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n462), .A2(new_n465), .B1(new_n208), .B2(G122), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n191), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n208), .A2(G122), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n468), .A2(new_n191), .A3(new_n469), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n459), .A2(new_n461), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n469), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(KEYINPUT14), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(G107), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n454), .A2(G134), .A3(new_n458), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G107), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n268), .A2(new_n269), .A3(new_n251), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n317), .B1(new_n479), .B2(new_n457), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n474), .A2(new_n475), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n375), .A2(new_n482), .A3(G953), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n471), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n471), .B2(new_n481), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n287), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT89), .B(new_n287), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n378), .A2(new_n445), .A3(new_n451), .A4(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n500));
  INV_X1    g314(.A(G131), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n320), .A2(G134), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n327), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n326), .A2(new_n276), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n265), .B1(new_n326), .B2(new_n329), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n265), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n330), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n323), .B2(new_n325), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n452), .A2(new_n453), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(new_n250), .B2(new_n252), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n511), .B1(new_n514), .B2(new_n344), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n273), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n517), .A3(KEYINPUT30), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n507), .A2(new_n518), .A3(new_n217), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n217), .A2(KEYINPUT71), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n215), .A2(new_n521), .A3(new_n216), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n509), .A2(new_n517), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n386), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT31), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n217), .B1(new_n505), .B2(new_n506), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n506), .B1(new_n334), .B2(new_n510), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n520), .A2(new_n522), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT28), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n528), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n507), .A2(new_n518), .A3(new_n217), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT31), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n523), .A4(new_n529), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n531), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT32), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT32), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n546), .A3(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n523), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n509), .A2(new_n517), .B1(new_n520), .B2(new_n522), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT28), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n537), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT29), .A4(new_n529), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n287), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n529), .B1(new_n534), .B2(new_n537), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n539), .A2(new_n523), .A3(new_n528), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G472), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n499), .B1(new_n548), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n542), .A2(new_n546), .A3(new_n543), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n546), .B1(new_n542), .B2(new_n543), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n499), .B(new_n558), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G110), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n270), .A2(KEYINPUT23), .A3(G119), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT23), .B1(new_n256), .B2(G119), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n256), .A2(G119), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n268), .A2(new_n269), .A3(new_n206), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(KEYINPUT24), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT24), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G110), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT74), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT74), .B1(new_n573), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n570), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n406), .A2(new_n408), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n397), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n405), .B2(G146), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT76), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n566), .A2(new_n569), .A3(new_n565), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n576), .A2(new_n577), .B1(new_n571), .B2(new_n568), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n583), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n581), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n581), .B(new_n597), .C1(new_n588), .C2(new_n589), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n482), .B1(G234), .B2(new_n287), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(G902), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n601), .B(KEYINPUT77), .Z(new_n602));
  INV_X1    g416(.A(new_n599), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(new_n287), .A3(new_n598), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(KEYINPUT25), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n596), .A2(new_n606), .A3(new_n287), .A4(new_n598), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n564), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n498), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n203), .ZN(G3));
  INV_X1    g427(.A(new_n310), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n302), .B2(new_n308), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n491), .A2(new_n287), .ZN(new_n616));
  INV_X1    g430(.A(new_n483), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n456), .A2(G134), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n454), .A2(new_n458), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n472), .A2(G107), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n466), .A2(new_n191), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n620), .A2(new_n460), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n480), .A2(new_n475), .A3(new_n478), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n476), .B1(new_n462), .B2(new_n465), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n466), .A2(new_n625), .A3(new_n191), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n617), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n471), .A2(new_n481), .A3(new_n483), .ZN(new_n629));
  AOI21_X1  g443(.A(G902), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n616), .B1(new_n630), .B2(new_n491), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT33), .B1(new_n484), .B2(new_n485), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n628), .A2(new_n633), .A3(new_n629), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n634), .A3(G478), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT90), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n631), .B2(new_n635), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n445), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n615), .A2(new_n451), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n376), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n354), .B2(new_n363), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n372), .B1(new_n643), .B2(new_n365), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n642), .B1(new_n644), .B2(new_n371), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n542), .A2(new_n287), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G472), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n544), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n649), .A3(new_n610), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT91), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT34), .B(G104), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  NAND3_X1  g468(.A1(new_n433), .A2(new_n439), .A3(KEYINPUT92), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT92), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(KEYINPUT20), .C1(new_n430), .C2(new_n432), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n492), .B1(new_n488), .B2(new_n489), .ZN(new_n659));
  INV_X1    g473(.A(new_n495), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n444), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n658), .A2(new_n661), .A3(new_n450), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n309), .A2(new_n662), .A3(new_n310), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT93), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT93), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n615), .A2(new_n665), .A3(new_n662), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n650), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT35), .B(G107), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  OAI21_X1  g483(.A(KEYINPUT94), .B1(new_n595), .B2(KEYINPUT36), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT94), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT36), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n593), .A2(new_n672), .A3(new_n673), .A4(new_n594), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n671), .B1(new_n670), .B2(new_n674), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n677), .B(new_n581), .C1(new_n589), .C2(new_n588), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n590), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n678), .A2(new_n680), .A3(new_n600), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n605), .B2(new_n607), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n440), .A2(new_n444), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n682), .A2(new_n683), .A3(new_n496), .A4(new_n450), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n378), .A2(new_n649), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT96), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n448), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n447), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n658), .A2(new_n661), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n681), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n608), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n694), .A2(new_n374), .A3(new_n376), .A4(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n311), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT97), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n564), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n615), .A2(new_n645), .A3(new_n696), .A4(new_n694), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT73), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n562), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT97), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XNOR2_X1  g521(.A(new_n692), .B(KEYINPUT39), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n377), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n309), .B(KEYINPUT38), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT40), .B1(new_n377), .B2(new_n709), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n549), .A2(new_n529), .A3(new_n550), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(G902), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n528), .B1(new_n539), .B2(new_n523), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n560), .B2(new_n561), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT98), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n723), .B(new_n720), .C1(new_n560), .C2(new_n561), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n683), .A2(new_n496), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(new_n310), .A3(new_n682), .A4(new_n727), .ZN(new_n728));
  OR3_X1    g542(.A1(new_n715), .A2(new_n716), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n716), .B1(new_n715), .B2(new_n728), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n251), .ZN(G45));
  AOI211_X1 g546(.A(new_n642), .B(new_n682), .C1(new_n644), .C2(new_n371), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n632), .A2(G478), .A3(new_n634), .ZN(new_n735));
  INV_X1    g549(.A(new_n616), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n486), .B2(G478), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT90), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n683), .A3(new_n692), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n734), .A2(new_n309), .A3(new_n741), .A4(new_n310), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n734), .B1(new_n615), .B2(new_n741), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n564), .B(new_n733), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  NOR2_X1   g559(.A1(new_n365), .A2(KEYINPUT101), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n643), .A2(new_n747), .ZN(new_n748));
  AOI211_X1 g562(.A(G902), .B(new_n746), .C1(new_n354), .C2(new_n363), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n748), .A2(new_n749), .A3(new_n642), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n703), .A2(new_n562), .A3(new_n610), .A4(new_n750), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(new_n641), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT41), .B(G113), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  AOI21_X1  g568(.A(new_n751), .B1(new_n666), .B2(new_n664), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT102), .B(G116), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G18));
  NAND3_X1  g571(.A1(new_n703), .A2(new_n562), .A3(new_n684), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n615), .A2(new_n750), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  NOR4_X1   g577(.A1(new_n748), .A2(new_n749), .A3(new_n450), .A4(new_n642), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n543), .B(KEYINPUT103), .Z(new_n765));
  NAND2_X1  g579(.A1(new_n531), .A2(new_n541), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n529), .B1(new_n551), .B2(new_n552), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n647), .A2(new_n608), .A3(new_n602), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n764), .A2(new_n770), .A3(new_n615), .A4(new_n727), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  INV_X1    g586(.A(new_n741), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n696), .A2(new_n647), .A3(new_n768), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n696), .A2(new_n647), .A3(KEYINPUT104), .A4(new_n768), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n761), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  NAND3_X1  g594(.A1(new_n302), .A2(new_n308), .A3(new_n310), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n377), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n609), .B1(new_n548), .B2(new_n558), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n564), .A2(new_n610), .A3(new_n741), .A4(new_n782), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n501), .ZN(G33));
  NOR2_X1   g604(.A1(new_n704), .A2(new_n609), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n694), .B(KEYINPUT106), .Z(new_n792));
  AND3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n782), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n317), .ZN(G36));
  NAND2_X1  g608(.A1(new_n445), .A2(new_n740), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT43), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n648), .A2(new_n696), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n781), .B(KEYINPUT107), .Z(new_n800));
  OAI21_X1  g614(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n368), .A2(new_n370), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT45), .ZN(new_n804));
  OAI21_X1  g618(.A(G469), .B1(new_n803), .B2(KEYINPUT45), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n373), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT46), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n806), .A2(new_n807), .B1(new_n365), .B2(new_n643), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n807), .B2(new_n806), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n376), .A3(new_n708), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NOR2_X1   g626(.A1(new_n773), .A2(new_n610), .ZN(new_n813));
  INV_X1    g627(.A(new_n781), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n704), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n376), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n818), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n815), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n391), .ZN(G42));
  NOR2_X1   g637(.A1(new_n748), .A2(new_n749), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT49), .Z(new_n825));
  NAND3_X1  g639(.A1(new_n610), .A2(new_n310), .A3(new_n376), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n825), .A2(new_n795), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n725), .ZN(new_n828));
  INV_X1    g642(.A(new_n713), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n642), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n819), .A2(new_n821), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n796), .A2(new_n691), .A3(new_n769), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n800), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n824), .A2(new_n376), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n614), .B1(KEYINPUT115), .B2(KEYINPUT50), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n829), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n776), .A2(new_n777), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n796), .A2(new_n691), .A3(new_n835), .A4(new_n781), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n840), .A2(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n835), .A2(new_n781), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n828), .A2(new_n845), .A3(new_n610), .A4(new_n447), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT116), .Z(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n445), .A3(new_n639), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n834), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n834), .A2(new_n844), .A3(KEYINPUT51), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n843), .A2(new_n783), .ZN(new_n853));
  NOR2_X1   g667(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n446), .B(G953), .C1(new_n833), .C2(new_n761), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n855), .B(new_n856), .C1(new_n853), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n640), .B2(new_n847), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n851), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  OAI221_X1 g675(.A(new_n771), .B1(new_n758), .B2(new_n760), .C1(new_n641), .C2(new_n751), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n861), .B1(new_n862), .B2(new_n755), .ZN(new_n863));
  INV_X1    g677(.A(new_n789), .ZN(new_n864));
  INV_X1    g678(.A(new_n748), .ZN(new_n865));
  INV_X1    g679(.A(new_n749), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n451), .A4(new_n376), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n769), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n614), .B(new_n726), .C1(new_n308), .C2(new_n302), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n759), .A2(new_n761), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n664), .A2(new_n666), .ZN(new_n871));
  INV_X1    g685(.A(new_n751), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n873), .A3(new_n752), .A4(KEYINPUT113), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n863), .A2(new_n864), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT114), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n863), .A2(new_n877), .A3(new_n864), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT109), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n640), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n445), .A2(new_n639), .A3(KEYINPUT109), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT110), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n445), .A2(new_n496), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n882), .A2(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n451), .A3(new_n615), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n445), .A2(new_n451), .A3(new_n496), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n311), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n650), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n685), .B1(new_n498), .B2(new_n611), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n778), .A2(new_n782), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n733), .A2(new_n703), .A3(new_n562), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n444), .A2(new_n692), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n658), .A2(new_n496), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n814), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n793), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(new_n899), .A3(KEYINPUT53), .ZN(new_n900));
  XNOR2_X1  g714(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n901));
  AOI211_X1 g715(.A(new_n693), .B(new_n681), .C1(new_n607), .C2(new_n605), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n725), .A2(new_n869), .A3(new_n645), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n779), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n743), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n615), .A2(new_n734), .A3(new_n741), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT111), .B1(new_n908), .B2(new_n706), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n374), .A2(new_n902), .A3(new_n376), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n722), .B2(new_n724), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n869), .A2(new_n911), .B1(new_n778), .B2(new_n761), .ZN(new_n912));
  AND4_X1   g726(.A1(KEYINPUT111), .A2(new_n706), .A3(new_n744), .A4(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n901), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n700), .A2(new_n705), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n742), .A2(new_n743), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n779), .B(new_n903), .C1(new_n916), .C2(new_n894), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n900), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n870), .A2(new_n873), .A3(new_n752), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n864), .A2(new_n892), .A3(new_n923), .A4(new_n899), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT111), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n915), .B2(new_n917), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n706), .A2(new_n912), .A3(KEYINPUT111), .A4(new_n744), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n926), .A2(KEYINPUT52), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT52), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT53), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n880), .A2(new_n921), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n892), .A2(new_n923), .A3(new_n864), .A4(new_n899), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n918), .B1(new_n909), .B2(new_n913), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n926), .A2(KEYINPUT52), .A3(new_n927), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n914), .A2(new_n920), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n924), .A2(new_n931), .ZN(new_n941));
  OAI221_X1 g755(.A(KEYINPUT54), .B1(new_n938), .B2(new_n931), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n860), .A2(new_n934), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT118), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n446), .A2(new_n280), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n943), .A2(new_n944), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n830), .B1(new_n947), .B2(new_n948), .ZN(G75));
  NOR2_X1   g763(.A1(new_n932), .A2(new_n287), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(G210), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n247), .B(new_n284), .ZN(new_n952));
  XOR2_X1   g766(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n951), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n280), .A2(G952), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(G51));
  AND3_X1   g774(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n899), .ZN(new_n961));
  INV_X1    g775(.A(new_n901), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n926), .B2(new_n927), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(new_n919), .ZN(new_n964));
  OAI22_X1  g778(.A1(new_n938), .A2(KEYINPUT53), .B1(new_n964), .B2(new_n879), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n933), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n372), .B(KEYINPUT57), .Z(new_n967));
  OAI21_X1  g781(.A(new_n364), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n804), .A2(new_n805), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n950), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n959), .B1(new_n968), .B2(new_n970), .ZN(G54));
  NAND3_X1  g785(.A1(new_n950), .A2(KEYINPUT58), .A3(G475), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(new_n430), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n430), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n959), .ZN(G60));
  NAND2_X1  g789(.A1(new_n934), .A2(new_n942), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n616), .B(KEYINPUT59), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n632), .A3(new_n634), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT121), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n632), .A2(new_n634), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n965), .A2(KEYINPUT54), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n934), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n980), .B1(new_n984), .B2(new_n959), .ZN(new_n985));
  INV_X1    g799(.A(new_n959), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT121), .B(new_n986), .C1(new_n966), .C2(new_n982), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n979), .A2(new_n985), .A3(new_n987), .ZN(G63));
  AND2_X1   g802(.A1(new_n678), .A2(new_n680), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n990));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n965), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n965), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT123), .B1(new_n932), .B2(new_n992), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n596), .A2(new_n598), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n965), .A2(new_n990), .A3(new_n993), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n996), .A2(new_n1000), .A3(new_n986), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n996), .A2(new_n1000), .A3(KEYINPUT61), .A4(new_n986), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(G66));
  INV_X1    g819(.A(new_n449), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n280), .B1(new_n1006), .B2(G224), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n892), .A2(new_n923), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n280), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n306), .B(new_n242), .C1(G898), .C2(new_n280), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(G69));
  OAI21_X1  g825(.A(new_n885), .B1(new_n882), .B2(new_n883), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n791), .A2(new_n710), .A3(new_n814), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n811), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT124), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT124), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n811), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n822), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n744), .A2(new_n779), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n706), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n731), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT62), .B1(new_n731), .B2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n280), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n507), .A2(new_n518), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(new_n426), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G900), .A2(G953), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n819), .A2(new_n821), .ZN(new_n1031));
  INV_X1    g845(.A(new_n815), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n864), .ZN(new_n1034));
  INV_X1    g848(.A(new_n793), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n869), .A2(new_n783), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n811), .B(new_n1035), .C1(new_n810), .C2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1034), .A2(new_n1020), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1030), .B1(new_n1038), .B2(new_n280), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT126), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1028), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1026), .B1(new_n1023), .B2(new_n280), .ZN(new_n1043));
  OAI21_X1  g857(.A(KEYINPUT126), .B1(new_n1043), .B2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(G227), .ZN(new_n1046));
  OAI21_X1  g860(.A(G953), .B1(new_n1046), .B2(new_n689), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1047), .B1(new_n1026), .B2(KEYINPUT125), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1042), .A2(new_n1048), .A3(new_n1044), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(G72));
  NAND2_X1  g866(.A1(G472), .A2(G902), .ZN(new_n1053));
  XOR2_X1   g867(.A(new_n1053), .B(KEYINPUT63), .Z(new_n1054));
  OAI21_X1  g868(.A(new_n1054), .B1(new_n1023), .B2(new_n1008), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n1055), .A2(new_n719), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1038), .A2(new_n923), .A3(new_n892), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n556), .B1(new_n1057), .B2(new_n1054), .ZN(new_n1058));
  INV_X1    g872(.A(new_n556), .ZN(new_n1059));
  INV_X1    g873(.A(new_n1054), .ZN(new_n1060));
  NOR3_X1   g874(.A1(new_n1059), .A2(new_n719), .A3(new_n1060), .ZN(new_n1061));
  XOR2_X1   g875(.A(new_n1061), .B(KEYINPUT127), .Z(new_n1062));
  OAI221_X1 g876(.A(new_n1062), .B1(new_n938), .B2(new_n931), .C1(new_n940), .C2(new_n941), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1063), .ZN(new_n1064));
  NOR4_X1   g878(.A1(new_n1056), .A2(new_n1058), .A3(new_n959), .A4(new_n1064), .ZN(G57));
endmodule


