//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n206));
  XNOR2_X1  g0006(.A(new_n205), .B(new_n206), .ZN(new_n207));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT65), .B(G238), .Z(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G58), .A2(G232), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n207), .B(new_n213), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g0043(.A(KEYINPUT68), .B1(new_n243), .B2(new_n210), .ZN(new_n244));
  INV_X1    g0044(.A(new_n210), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT68), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n244), .A2(new_n247), .A3(G274), .A4(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n250), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n244), .A2(new_n252), .A3(new_n247), .A4(G232), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G87), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT75), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  MUX2_X1   g0059(.A(G223), .B(G226), .S(G1698), .Z(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n243), .A2(new_n210), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n251), .B(new_n253), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G190), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(G200), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n210), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT7), .B1(new_n259), .B2(G20), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n211), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n272), .A2(G68), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(G58), .B(G68), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n279), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT16), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT16), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(new_n284), .A3(new_n281), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n271), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G1), .B2(new_n211), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n270), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n290), .A2(new_n294), .B1(new_n293), .B2(new_n287), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n286), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT76), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT17), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n268), .A2(new_n297), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n285), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n284), .B1(new_n278), .B2(new_n281), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n270), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n305), .A2(new_n266), .A3(new_n295), .A4(new_n267), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(new_n299), .A3(new_n300), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n264), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n260), .A2(new_n259), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n262), .B1(new_n312), .B2(new_n256), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n251), .A4(new_n253), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT18), .B1(new_n297), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n305), .A2(new_n295), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT18), .ZN(new_n319));
  INV_X1    g0119(.A(new_n316), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n308), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n211), .A2(G33), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n288), .ZN(new_n326));
  INV_X1    g0126(.A(G50), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n215), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n270), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n292), .A2(G50), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n270), .B1(new_n291), .B2(G20), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(G50), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n339), .B(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n244), .A2(new_n247), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G226), .A3(new_n252), .ZN(new_n343));
  INV_X1    g0143(.A(G1698), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n257), .B2(new_n258), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G223), .ZN(new_n346));
  INV_X1    g0146(.A(G77), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n259), .ZN(new_n348));
  AOI21_X1  g0148(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(G222), .B2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n251), .B(new_n343), .C1(new_n350), .C2(new_n263), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n265), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G200), .B2(new_n351), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT10), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n341), .A2(new_n353), .B1(KEYINPUT72), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(KEYINPUT72), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n341), .A2(new_n359), .A3(KEYINPUT10), .A4(new_n353), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n339), .B1(new_n309), .B2(new_n351), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G179), .B2(new_n351), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT71), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n287), .B(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n366), .A2(new_n280), .ZN(new_n367));
  INV_X1    g0167(.A(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT15), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT15), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n373), .A2(new_n324), .B1(new_n211), .B2(new_n347), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n270), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n292), .A2(G77), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n335), .B2(G77), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n342), .A2(G244), .A3(new_n252), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(new_n251), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n259), .A2(G232), .A3(new_n344), .ZN(new_n381));
  INV_X1    g0181(.A(G107), .ZN(new_n382));
  INV_X1    g0182(.A(new_n345), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n381), .B1(new_n382), .B2(new_n259), .C1(new_n383), .C2(new_n214), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n262), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n378), .B1(G200), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(G190), .A3(new_n385), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n386), .A2(new_n309), .B1(new_n375), .B2(new_n377), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n380), .A2(new_n314), .A3(new_n385), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n387), .A2(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n349), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n263), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n244), .A2(new_n252), .A3(new_n247), .A4(G238), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n251), .ZN(new_n396));
  OR3_X1    g0196(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT13), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT13), .B1(new_n394), .B2(new_n396), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G169), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n398), .A2(new_n402), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n403), .A2(G179), .A3(new_n404), .A4(new_n397), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(new_n406), .A3(G169), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n325), .A2(G77), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n280), .A2(G50), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n211), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(KEYINPUT74), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(KEYINPUT74), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n270), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT11), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  OR3_X1    g0217(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT12), .B1(new_n292), .B2(G68), .ZN(new_n419));
  AOI22_X1  g0219(.A1(G68), .A2(new_n335), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n408), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(G200), .B2(new_n399), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n403), .A2(new_n404), .A3(new_n397), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n265), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AND4_X1   g0226(.A1(new_n323), .A2(new_n364), .A3(new_n391), .A4(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n345), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n428));
  OAI211_X1 g0228(.A(G244), .B(new_n344), .C1(new_n273), .C2(new_n274), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT80), .B1(new_n429), .B2(KEYINPUT79), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT4), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n429), .B2(KEYINPUT80), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(KEYINPUT80), .B(new_n431), .C1(new_n429), .C2(KEYINPUT79), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n262), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n291), .A2(G45), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT5), .A2(G41), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n441), .A2(G257), .A3(new_n244), .A4(new_n247), .ZN(new_n442));
  INV_X1    g0242(.A(new_n440), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n443), .B2(new_n438), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n444), .A2(G274), .A3(new_n244), .A4(new_n247), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n435), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n265), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n429), .A2(KEYINPUT79), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT80), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT4), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n428), .C1(new_n430), .C2(new_n432), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n446), .B1(new_n453), .B2(new_n262), .ZN(new_n454));
  INV_X1    g0254(.A(G200), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n272), .A2(G107), .A3(new_n277), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT78), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT6), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n382), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n382), .A2(KEYINPUT6), .A3(G97), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n211), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n280), .A2(G77), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT77), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT78), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n272), .A2(new_n277), .A3(new_n469), .A4(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n270), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n292), .A2(G97), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n291), .A2(G33), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n294), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n476), .B2(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n449), .A2(new_n456), .A3(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n314), .B(new_n446), .C1(new_n453), .C2(new_n262), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n309), .B1(new_n435), .B2(new_n447), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT81), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT81), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n478), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n479), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT83), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n345), .A2(new_n487), .A3(G264), .ZN(new_n488));
  OAI211_X1 g0288(.A(G264), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n349), .A2(G257), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n275), .A2(G303), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n262), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n441), .A2(G270), .A3(new_n244), .A4(new_n247), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n445), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(G20), .B1(G33), .B2(G283), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G33), .B2(new_n460), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G20), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n270), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n476), .A2(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n293), .A2(new_n501), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n498), .A2(new_n508), .A3(KEYINPUT21), .A4(G169), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n262), .B2(new_n493), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n510), .A3(G179), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n503), .B(KEYINPUT20), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n507), .B1(new_n475), .B2(new_n501), .ZN(new_n515));
  OAI21_X1  g0315(.A(G169), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n494), .A2(new_n497), .A3(G190), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n510), .C2(new_n455), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n512), .A2(KEYINPUT84), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n517), .A3(new_n509), .A4(new_n511), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT84), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n259), .A2(new_n211), .A3(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n529), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n259), .A2(new_n211), .A3(G87), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(new_n382), .A3(G20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT87), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n527), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT87), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n538), .B(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(new_n526), .A3(new_n530), .A4(new_n532), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n271), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n382), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT25), .B1(new_n293), .B2(new_n382), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n475), .A2(new_n382), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G250), .B(new_n344), .C1(new_n273), .C2(new_n274), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G294), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n262), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n441), .A2(G264), .A3(new_n244), .A4(new_n247), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n445), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n309), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G179), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT82), .ZN(new_n559));
  NAND3_X1  g0359(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n211), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n462), .A2(new_n368), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n211), .B(G68), .C1(new_n273), .C2(new_n274), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n324), .B2(new_n460), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n270), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n372), .A2(new_n292), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n559), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI211_X1 g0372(.A(KEYINPUT82), .B(new_n569), .C1(new_n567), .C2(new_n270), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n572), .A2(new_n574), .B1(new_n372), .B2(new_n476), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n244), .A2(new_n247), .A3(G274), .A4(new_n437), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n244), .A2(new_n247), .A3(G250), .A4(new_n436), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n345), .A2(G244), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n259), .A2(G238), .A3(new_n344), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G116), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n262), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(new_n584), .A3(new_n314), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n578), .B1(new_n262), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(G169), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n584), .A3(G190), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n586), .B2(new_n455), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n476), .A2(G87), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n571), .B2(new_n573), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n575), .A2(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n555), .A2(G200), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n553), .A2(G190), .A3(new_n445), .A4(new_n554), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n544), .A2(new_n595), .A3(new_n547), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n558), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n427), .A2(new_n486), .A3(new_n525), .A4(new_n597), .ZN(G372));
  NAND2_X1  g0398(.A1(new_n389), .A2(new_n390), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n425), .A2(new_n600), .B1(new_n408), .B2(new_n421), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n308), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n358), .B(new_n360), .C1(new_n602), .C2(new_n322), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n362), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT91), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n483), .A2(new_n485), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT88), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n591), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(KEYINPUT88), .B(new_n590), .C1(new_n571), .C2(new_n573), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n589), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n575), .A2(new_n587), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n611), .A2(new_n596), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT89), .ZN(new_n614));
  OR3_X1    g0414(.A1(new_n449), .A2(new_n456), .A3(new_n478), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n607), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n512), .A2(new_n517), .ZN(new_n617));
  INV_X1    g0417(.A(new_n558), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n614), .B1(new_n486), .B2(new_n613), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT26), .B1(new_n607), .B2(new_n592), .ZN(new_n623));
  INV_X1    g0423(.A(new_n612), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n611), .A2(new_n612), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n435), .A2(G179), .A3(new_n447), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(KEYINPUT90), .C1(new_n309), .C2(new_n454), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n472), .A2(new_n477), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n309), .B2(new_n454), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n625), .A2(new_n626), .A3(new_n628), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n623), .A2(new_n624), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n427), .B1(new_n622), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n606), .A2(new_n635), .ZN(G369));
  NAND3_X1  g0436(.A1(new_n291), .A2(new_n211), .A3(G13), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G213), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(G343), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n617), .A2(new_n519), .A3(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n521), .A2(new_n524), .B1(new_n508), .B2(new_n642), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n618), .A2(new_n642), .ZN(new_n647));
  INV_X1    g0447(.A(new_n596), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n642), .B1(new_n544), .B2(new_n547), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n558), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G330), .ZN(new_n652));
  OR3_X1    g0452(.A1(new_n646), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT92), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n617), .A2(new_n642), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  OR3_X1    g0458(.A1(new_n657), .A2(new_n658), .A3(new_n647), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n657), .B2(new_n647), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n655), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n204), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n663), .A2(KEYINPUT94), .A3(G41), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT94), .B1(new_n663), .B2(G41), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n562), .A2(G116), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n666), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n209), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT28), .Z(new_n671));
  INV_X1    g0471(.A(new_n485), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n484), .B1(new_n630), .B2(new_n478), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n592), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n626), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n632), .A2(new_n628), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n611), .A2(new_n612), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n679), .A3(new_n624), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT98), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n619), .A2(new_n486), .A3(new_n613), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n680), .B2(new_n681), .ZN(new_n684));
  OAI211_X1 g0484(.A(KEYINPUT29), .B(new_n643), .C1(new_n682), .C2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n615), .B1(new_n672), .B2(new_n673), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n625), .A2(new_n648), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT89), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n616), .A3(new_n619), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n626), .B1(new_n674), .B2(new_n675), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n633), .A2(new_n624), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n642), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n685), .B1(KEYINPUT29), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n579), .A2(new_n584), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n498), .A2(new_n314), .A3(new_n696), .A4(new_n555), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n454), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n553), .A2(new_n554), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n510), .A2(G179), .A3(new_n586), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT30), .B1(new_n700), .B2(new_n448), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n494), .A2(new_n497), .A3(G179), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n579), .A2(new_n584), .A3(new_n553), .A4(new_n554), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n454), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n698), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT96), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n642), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI211_X1 g0509(.A(KEYINPUT96), .B(new_n698), .C1(new_n701), .C2(new_n706), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n695), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n525), .A2(new_n486), .A3(new_n597), .A4(new_n643), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n701), .A2(new_n706), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n697), .A2(new_n454), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n643), .A2(new_n695), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n716), .A2(KEYINPUT95), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT95), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n712), .A2(new_n713), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n711), .A2(KEYINPUT97), .ZN(new_n722));
  OAI21_X1  g0522(.A(G330), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n694), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n671), .B1(new_n724), .B2(G1), .ZN(G364));
  INV_X1    g0525(.A(G13), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n291), .B1(new_n727), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n669), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT100), .ZN(new_n732));
  OAI21_X1  g0532(.A(G20), .B1(new_n732), .B2(G169), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n309), .A2(KEYINPUT100), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n245), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n211), .A2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(G179), .A3(new_n455), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n275), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n211), .A2(new_n265), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n314), .A2(new_n455), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G326), .ZN(new_n750));
  INV_X1    g0550(.A(new_n746), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(new_n455), .A3(G179), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n211), .B1(new_n756), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n745), .B(new_n755), .C1(G294), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n314), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n746), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n740), .A2(new_n760), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n740), .A2(new_n756), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G329), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n747), .A2(new_n740), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT102), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT103), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n759), .B(new_n768), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT104), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(G159), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n753), .A2(new_n368), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n757), .A2(new_n460), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n781), .A2(new_n782), .A3(new_n275), .A4(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n748), .A2(new_n327), .B1(new_n761), .B2(new_n328), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n743), .A2(new_n382), .B1(new_n763), .B2(new_n347), .ZN(new_n786));
  INV_X1    g0586(.A(new_n774), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n785), .B(new_n786), .C1(G68), .C2(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n777), .A2(new_n778), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n739), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n738), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n259), .A2(new_n204), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G355), .B1(new_n501), .B2(new_n663), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n237), .A2(new_n249), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n663), .A2(new_n259), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n208), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n731), .B(new_n790), .C1(new_n794), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n646), .ZN(new_n803));
  INV_X1    g0603(.A(new_n793), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT105), .Z(new_n806));
  OAI21_X1  g0606(.A(new_n731), .B1(new_n646), .B2(new_n652), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n652), .B2(new_n646), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  OAI21_X1  g0610(.A(KEYINPUT108), .B1(new_n599), .B2(new_n643), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT108), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n389), .A2(new_n812), .A3(new_n390), .A4(new_n642), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n378), .A2(new_n642), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n811), .A2(new_n813), .B1(new_n391), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n693), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n730), .B1(new_n817), .B2(new_n723), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n723), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n738), .A2(new_n791), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n731), .B1(new_n820), .B2(new_n347), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n259), .B1(new_n753), .B2(new_n327), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n743), .A2(new_n215), .B1(new_n766), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n328), .B2(new_n757), .ZN(new_n826));
  INV_X1    g0626(.A(new_n761), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G137), .A2(new_n749), .B1(new_n827), .B2(G143), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n763), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G150), .B2(new_n787), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n826), .B1(KEYINPUT34), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n748), .A2(new_n754), .B1(new_n763), .B2(new_n501), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n787), .B2(G283), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT106), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n752), .A2(G107), .B1(G294), .B2(new_n827), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n764), .B2(new_n766), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n743), .A2(new_n368), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n838), .A2(new_n259), .A3(new_n783), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n832), .A2(new_n833), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n739), .B1(new_n841), .B2(KEYINPUT107), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n841), .A2(KEYINPUT107), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n821), .B1(new_n816), .B2(new_n792), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n819), .A2(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n727), .A2(new_n291), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n716), .A2(KEYINPUT96), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n707), .A2(new_n708), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(KEYINPUT31), .A3(new_n642), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n711), .A2(new_n851), .A3(new_n713), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n421), .A2(new_n642), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n422), .A2(new_n425), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n408), .A2(new_n421), .A3(new_n642), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n815), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n640), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n286), .B2(new_n296), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n308), .B2(new_n322), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n318), .A2(new_n320), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n306), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n306), .A3(new_n865), .A4(new_n859), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n861), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n848), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n869), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n861), .A2(new_n867), .A3(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n852), .A4(new_n856), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT110), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n427), .A2(new_n852), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(G330), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n854), .A2(new_n855), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n599), .A2(new_n642), .ZN(new_n883));
  AOI211_X1 g0683(.A(KEYINPUT109), .B(new_n883), .C1(new_n693), .C2(new_n816), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT109), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n643), .B(new_n816), .C1(new_n622), .C2(new_n634), .ZN(new_n886));
  INV_X1    g0686(.A(new_n883), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n874), .B(new_n882), .C1(new_n884), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n874), .B(KEYINPUT39), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n422), .A2(new_n642), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n890), .A2(new_n891), .B1(new_n322), .B2(new_n640), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n427), .B(new_n685), .C1(KEYINPUT29), .C2(new_n693), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n606), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n847), .B1(new_n881), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n881), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n463), .A2(new_n464), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(KEYINPUT35), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(G116), .A3(new_n212), .A4(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT36), .ZN(new_n903));
  OAI21_X1  g0703(.A(G77), .B1(new_n328), .B2(new_n215), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n904), .A2(new_n208), .B1(G50), .B2(new_n215), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(G1), .A3(new_n726), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n903), .A3(new_n906), .ZN(G367));
  NAND3_X1  g0707(.A1(new_n609), .A2(new_n610), .A3(new_n642), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n624), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n625), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n793), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n232), .A2(new_n799), .B1(new_n663), .B2(new_n372), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n731), .B1(new_n794), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(G150), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n753), .A2(new_n328), .B1(new_n761), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n275), .B(new_n915), .C1(G143), .C2(new_n749), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n758), .A2(G68), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n787), .A2(G159), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n743), .A2(new_n347), .B1(new_n763), .B2(new_n327), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G137), .B2(new_n767), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT112), .B1(new_n753), .B2(new_n501), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT46), .Z(new_n923));
  INV_X1    g0723(.A(G294), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n924), .B2(new_n774), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n259), .B1(new_n742), .B2(G97), .ZN(new_n926));
  INV_X1    g0726(.A(new_n763), .ZN(new_n927));
  AOI22_X1  g0727(.A1(G303), .A2(new_n827), .B1(new_n927), .B2(G283), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n749), .A2(G311), .B1(new_n767), .B2(G317), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n758), .A2(G107), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n926), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n921), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n738), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n911), .B(new_n913), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n486), .B1(new_n629), .B2(new_n643), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n632), .A2(new_n628), .A3(new_n642), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n659), .A2(new_n660), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT44), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n661), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT45), .B1(new_n661), .B2(new_n940), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(new_n655), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n646), .A2(new_n652), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(KEYINPUT111), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n651), .B(new_n656), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n950), .B(KEYINPUT111), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n724), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n724), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n666), .B(KEYINPUT41), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n729), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n657), .A2(new_n940), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n940), .A2(new_n558), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n642), .B1(new_n963), .B2(new_n607), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT43), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n962), .A2(new_n964), .B1(new_n965), .B2(new_n910), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n910), .A2(new_n965), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n655), .A2(new_n941), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n937), .B1(new_n960), .B2(new_n970), .ZN(G387));
  NOR2_X1   g0771(.A1(new_n763), .A2(new_n215), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n753), .A2(new_n347), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G159), .C2(new_n749), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n373), .A2(new_n757), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n761), .A2(new_n327), .B1(new_n766), .B2(new_n914), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n275), .B(new_n977), .C1(G97), .C2(new_n742), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n787), .A2(new_n288), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n259), .B1(new_n767), .B2(G326), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n752), .A2(G294), .B1(G283), .B2(new_n758), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT115), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G317), .A2(new_n827), .B1(new_n927), .B2(G303), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n762), .B2(new_n748), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G311), .B2(new_n787), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n983), .B1(new_n986), .B2(KEYINPUT48), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT48), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT49), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n981), .B1(new_n501), .B2(new_n743), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n980), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n738), .ZN(new_n993));
  INV_X1    g0793(.A(new_n229), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n799), .B1(new_n994), .B2(new_n249), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n366), .A2(new_n327), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT114), .Z(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n667), .B(new_n249), .C1(new_n215), .C2(new_n347), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n997), .B2(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n995), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n796), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n667), .B1(G107), .B2(new_n204), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n794), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n993), .A2(new_n730), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n651), .B2(new_n793), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n955), .B2(new_n729), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n956), .A2(new_n669), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n724), .A2(new_n955), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(G393));
  NAND2_X1  g0810(.A1(new_n949), .A2(new_n956), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n956), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n666), .B1(new_n948), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n767), .A2(G143), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n753), .B2(new_n215), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n757), .A2(new_n347), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1016), .A2(new_n839), .A3(new_n1017), .A4(new_n275), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n748), .A2(new_n914), .B1(new_n761), .B2(new_n829), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT51), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n787), .A2(G50), .B1(new_n366), .B2(new_n927), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n753), .A2(new_n744), .B1(new_n766), .B2(new_n762), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G294), .B2(new_n927), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n275), .B1(new_n743), .B2(new_n382), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G116), .B2(new_n758), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(new_n754), .C2(new_n774), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G317), .A2(new_n749), .B1(new_n827), .B2(G311), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT52), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1022), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1030), .A2(new_n738), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n240), .A2(new_n799), .B1(G97), .B2(new_n663), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n731), .B(new_n1031), .C1(new_n794), .C2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n940), .B2(new_n804), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n949), .B2(new_n728), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1014), .A2(new_n1035), .ZN(G390));
  INV_X1    g0836(.A(new_n882), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n723), .B2(new_n815), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n852), .A2(new_n856), .A3(G330), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n642), .B(new_n815), .C1(new_n689), .C2(new_n692), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT109), .B1(new_n1041), .B2(new_n883), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n886), .A2(new_n885), .A3(new_n887), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n643), .B1(new_n716), .B2(KEYINPUT96), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT31), .B1(new_n1046), .B2(new_n850), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT97), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1049), .A2(new_n712), .A3(new_n713), .A4(new_n720), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1050), .A2(new_n882), .A3(G330), .A4(new_n816), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n852), .A2(G330), .A3(new_n816), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n1037), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n643), .B(new_n816), .C1(new_n682), .C2(new_n684), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n887), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1045), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n427), .A2(G330), .A3(new_n852), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n606), .A2(new_n894), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT116), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n882), .B1(new_n884), .B2(new_n888), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n891), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n890), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n870), .B(new_n891), .C1(new_n1056), .C2(new_n882), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1051), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n890), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n891), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n874), .B(new_n1065), .C1(new_n1057), .C2(new_n1037), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1039), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT116), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1044), .A2(new_n1040), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n1061), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1039), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1072), .A2(new_n1073), .A3(new_n1051), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1075), .A2(new_n669), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n729), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n757), .A2(new_n829), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n753), .A2(new_n914), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1087));
  OAI221_X1 g0887(.A(new_n259), .B1(new_n823), .B2(new_n761), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(KEYINPUT54), .B(G143), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n787), .A2(G137), .B1(new_n927), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(G125), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n743), .A2(new_n327), .B1(new_n766), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G128), .B2(new_n749), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1089), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n774), .A2(new_n382), .B1(new_n460), .B2(new_n763), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT119), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n742), .A2(G68), .B1(new_n827), .B2(G116), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n749), .A2(G283), .B1(new_n767), .B2(G294), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n782), .A2(new_n259), .A3(new_n1017), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1098), .A2(new_n1099), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n738), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n731), .B1(new_n820), .B2(new_n287), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n890), .C2(new_n792), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1084), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1083), .A2(new_n1112), .ZN(G378));
  NAND3_X1  g0913(.A1(new_n1080), .A2(new_n1081), .A3(new_n1059), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1062), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n871), .A2(new_n875), .A3(G330), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n858), .B1(new_n337), .B2(new_n338), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n363), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1121));
  NAND4_X1  g0921(.A1(new_n358), .A2(new_n360), .A3(new_n362), .A4(new_n1118), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1116), .B(KEYINPUT123), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1116), .A2(KEYINPUT123), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT123), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n871), .A2(new_n875), .A3(new_n1128), .A4(G330), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1125), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(new_n893), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1115), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n889), .A3(new_n892), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n893), .B(new_n1125), .C1(new_n1126), .C2(new_n1130), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n666), .B1(new_n1115), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1127), .A2(new_n791), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G33), .B(G41), .C1(new_n742), .C2(G159), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n752), .A2(new_n1091), .B1(G137), .B2(new_n927), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n761), .C1(new_n774), .C2(new_n823), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n748), .A2(new_n1095), .B1(new_n757), .B2(new_n914), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT120), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1144), .B(new_n1152), .C1(G124), .C2(new_n767), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G116), .A2(new_n749), .B1(new_n827), .B2(G107), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n744), .B2(new_n766), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n743), .A2(new_n328), .B1(new_n373), .B2(new_n763), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1156), .A2(new_n973), .A3(G41), .A4(new_n259), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n917), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1155), .B(new_n1158), .C1(G97), .C2(new_n787), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT58), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(KEYINPUT58), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n327), .B1(new_n273), .B2(G41), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n738), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n731), .B1(new_n820), .B2(new_n327), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1142), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1132), .B2(new_n728), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1141), .A2(new_n1169), .ZN(G375));
  NAND2_X1  g0970(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1077), .A2(new_n1061), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n959), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n748), .A2(new_n924), .B1(new_n763), .B2(new_n382), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n787), .B2(G116), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT124), .Z(new_n1176));
  AOI22_X1  g0976(.A1(G283), .A2(new_n827), .B1(new_n767), .B2(G303), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n460), .B2(new_n753), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n275), .B1(new_n743), .B2(new_n347), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n975), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n758), .A2(G50), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n753), .A2(new_n829), .B1(new_n766), .B2(new_n1146), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n275), .B(new_n1182), .C1(G58), .C2(new_n742), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n787), .A2(new_n1091), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n748), .A2(new_n823), .B1(new_n763), .B2(new_n914), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G137), .B2(new_n827), .ZN(new_n1186));
  AND4_X1   g0986(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .A4(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n738), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n731), .B1(new_n820), .B2(new_n215), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n882), .C2(new_n792), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1077), .B2(new_n728), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1173), .A2(new_n1192), .ZN(G381));
  NOR2_X1   g0993(.A1(new_n1014), .A2(new_n1035), .ZN(new_n1194));
  INV_X1    g0994(.A(G384), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1196), .A2(G396), .A3(G393), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT125), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1083), .A2(new_n1198), .A3(new_n1112), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1083), .B2(new_n1112), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1169), .A3(new_n1141), .ZN(new_n1202));
  OR4_X1    g1002(.A1(G387), .A2(new_n1197), .A3(new_n1202), .A4(G381), .ZN(G407));
  OAI211_X1 g1003(.A(G407), .B(G213), .C1(G343), .C2(new_n1202), .ZN(G409));
  OAI211_X1 g1004(.A(G390), .B(new_n937), .C1(new_n960), .C2(new_n970), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(G393), .B(new_n809), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(G387), .A2(new_n1194), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT61), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n641), .A2(G213), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(G2897), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n1061), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n669), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1171), .A2(KEYINPUT60), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1172), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1195), .B1(new_n1218), .B2(new_n1191), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1217), .A2(new_n1172), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G384), .B(new_n1192), .C1(new_n1220), .C2(new_n1216), .ZN(new_n1221));
  AOI211_X1 g1021(.A(KEYINPUT127), .B(new_n1214), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT127), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G2897), .B(new_n1213), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1132), .B1(new_n1062), .B2(new_n1114), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1168), .B1(new_n1228), .B2(new_n959), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1199), .A2(new_n1229), .A3(new_n1200), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1115), .A2(new_n1139), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n669), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT57), .B1(new_n1115), .B2(new_n1133), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1169), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT126), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1141), .A2(new_n1236), .A3(G378), .A4(new_n1169), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1230), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1227), .B1(new_n1238), .B2(new_n1213), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1238), .A2(new_n1213), .A3(new_n1223), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT62), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1211), .B(new_n1239), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1230), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1223), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1212), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(KEYINPUT62), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1210), .B1(new_n1242), .B2(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1239), .A2(new_n1211), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1240), .A2(KEYINPUT63), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n1255), .ZN(G405));
  NAND2_X1  g1056(.A1(G375), .A2(new_n1201), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1243), .A2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(new_n1223), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(new_n1251), .ZN(G402));
endmodule


