//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR3_X1   g035(.A1(new_n459), .A2(new_n460), .A3(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT66), .B1(new_n462), .B2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G101), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G137), .A3(new_n462), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n477));
  OR3_X1    g052(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n468), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n468), .A2(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n480), .B(new_n484), .C1(G136), .C2(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(KEYINPUT68), .A2(KEYINPUT4), .A3(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n466), .B2(new_n467), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n462), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n466), .B2(new_n467), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n462), .C1(new_n471), .C2(new_n472), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT68), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n492), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT69), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(new_n509), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n516), .A2(new_n506), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n513), .A2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n517), .A2(G89), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n514), .A2(new_n512), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n519), .A2(G63), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(new_n525), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n517), .A2(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n524), .A2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n506), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(G43), .A2(new_n524), .B1(new_n517), .B2(G81), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n516), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(KEYINPUT70), .B(new_n538), .C1(new_n516), .C2(new_n539), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G651), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND4_X1  g126(.A1(new_n508), .A2(G53), .A3(G543), .A4(new_n509), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(KEYINPUT71), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n552), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n516), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n517), .A2(G91), .B1(new_n558), .B2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G299));
  NAND3_X1  g135(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(G301));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND3_X1  g137(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT72), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n515), .A2(G74), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n517), .A2(G87), .B1(G651), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(new_n524), .A2(G48), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n517), .A2(G86), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n506), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT73), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(new_n517), .A2(G85), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n524), .A2(G47), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n506), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n517), .A2(G92), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT75), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n516), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n524), .A2(G54), .B1(new_n588), .B2(G651), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n580), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n580), .B1(new_n591), .B2(G868), .ZN(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(G299), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n591), .B1(new_n598), .B2(G860), .ZN(G148));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n545), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n590), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g179(.A1(new_n461), .A2(new_n463), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n468), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT13), .Z(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(G2100), .ZN(new_n611));
  AOI22_X1  g186(.A1(G123), .A2(new_n482), .B1(new_n486), .B2(G135), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(G111), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(KEYINPUT77), .B1(new_n614), .B2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT77), .B2(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n610), .A2(new_n611), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT78), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n622), .B2(new_n623), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT79), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n632), .B(new_n633), .Z(new_n634));
  OR2_X1    g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n636), .A3(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n639), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  OAI221_X1 g221(.A(new_n641), .B1(new_n640), .B2(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n641), .A2(new_n643), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(new_n618), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT20), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G1986), .Z(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n666), .B(new_n667), .ZN(new_n673));
  INV_X1    g248(.A(new_n671), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NOR2_X1   g252(.A1(G171), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G5), .B2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(G1961), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT31), .B(G11), .Z(new_n682));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(G28), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n685), .A2(new_n686), .B1(new_n684), .B2(G28), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n682), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G168), .A2(new_n677), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n677), .B2(G21), .ZN(new_n691));
  INV_X1    g266(.A(G1966), .ZN(new_n692));
  OAI221_X1 g267(.A(new_n689), .B1(new_n683), .B2(new_n617), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n681), .B(new_n693), .C1(new_n692), .C2(new_n691), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n683), .A2(G35), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n683), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT29), .Z(new_n698));
  INV_X1    g273(.A(G2090), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G27), .A2(G29), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G164), .B2(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G2078), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n683), .A2(G32), .ZN(new_n704));
  AOI22_X1  g279(.A1(G129), .A2(new_n482), .B1(new_n605), .B2(G105), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n486), .A2(G141), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n683), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT27), .B(G1996), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G2078), .ZN(new_n714));
  INV_X1    g289(.A(new_n702), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n683), .A2(G33), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT25), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(new_n462), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n719), .B(new_n721), .C1(G139), .C2(new_n486), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n717), .B1(new_n722), .B2(new_n683), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2072), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  OAI21_X1  g300(.A(G29), .B1(new_n470), .B2(new_n475), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n724), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n700), .A2(new_n703), .A3(new_n716), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n679), .A2(new_n680), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(G2084), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT88), .Z(new_n737));
  OAI211_X1 g312(.A(new_n735), .B(new_n737), .C1(new_n698), .C2(new_n699), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n677), .A2(G20), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1956), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n734), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n677), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n546), .B2(new_n677), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT86), .B(G1341), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(G104), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n751));
  INV_X1    g326(.A(G140), .ZN(new_n752));
  INV_X1    g327(.A(G128), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n751), .B1(new_n485), .B2(new_n752), .C1(new_n753), .C2(new_n481), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n683), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n677), .A2(G4), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n591), .B2(new_n677), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n759), .B1(new_n761), .B2(G1348), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n749), .B(new_n762), .C1(G1348), .C2(new_n761), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT87), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n695), .A2(new_n745), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n677), .A2(G23), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G288), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT84), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT33), .B(G1976), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n677), .A2(G22), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G166), .B2(new_n677), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1971), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT32), .B(G1981), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n677), .A2(G6), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n573), .B2(new_n677), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT34), .B1(new_n771), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n486), .A2(G131), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n482), .A2(G119), .ZN(new_n782));
  NOR2_X1   g357(.A1(G95), .A2(G2105), .ZN(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n683), .A2(G25), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT81), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT82), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n677), .A2(G24), .ZN(new_n793));
  INV_X1    g368(.A(G290), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n677), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT83), .Z(new_n796));
  OAI21_X1  g371(.A(new_n792), .B1(G1986), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G1986), .B2(new_n796), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n780), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n771), .A2(new_n779), .A3(KEYINPUT34), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n766), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n804), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n806), .A2(KEYINPUT36), .A3(new_n802), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n765), .B1(new_n805), .B2(new_n807), .ZN(G311));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  INV_X1    g384(.A(new_n765), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(G150));
  NAND2_X1  g386(.A1(new_n517), .A2(G93), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n524), .A2(G55), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(new_n506), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT92), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n545), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n546), .A2(new_n817), .A3(new_n816), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT38), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n591), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT93), .B(G860), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n816), .A2(new_n828), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  NAND2_X1  g408(.A1(new_n482), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G142), .B2(new_n486), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n785), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n710), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n754), .B(new_n501), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n722), .ZN(new_n842));
  INV_X1    g417(.A(new_n608), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n840), .A2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n617), .B(G160), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G162), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  INV_X1    g426(.A(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g430(.A(new_n573), .B(G303), .ZN(new_n856));
  NAND2_X1  g431(.A1(G288), .A2(G290), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(G288), .A2(G290), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT94), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n856), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n858), .A2(KEYINPUT94), .A3(new_n859), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n573), .B(G166), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT42), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n823), .B(new_n602), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n590), .A2(new_n595), .ZN(new_n873));
  NAND4_X1  g448(.A1(G299), .A2(new_n584), .A3(new_n585), .A4(new_n589), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n875), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n879), .B2(new_n872), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT42), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n871), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n871), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G868), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n816), .A2(G868), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G295));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n885), .B2(new_n887), .ZN(new_n890));
  AOI211_X1 g465(.A(KEYINPUT96), .B(new_n886), .C1(new_n884), .C2(G868), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n821), .A2(new_n822), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n821), .B2(new_n822), .ZN(new_n896));
  OR3_X1    g471(.A1(G171), .A2(KEYINPUT97), .A3(G286), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT97), .B1(G171), .B2(G286), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT98), .B1(G168), .B2(G301), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n901));
  NAND3_X1  g476(.A1(G171), .A2(new_n901), .A3(G286), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n895), .A2(new_n896), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n823), .A2(KEYINPUT99), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n897), .A2(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n821), .A2(new_n822), .A3(new_n894), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n904), .A2(new_n879), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n876), .B1(new_n904), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n911), .B2(new_n868), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(new_n879), .A3(new_n908), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n910), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n904), .A2(new_n879), .A3(new_n908), .A4(KEYINPUT102), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n864), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT101), .B1(new_n864), .B2(new_n867), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n918), .A2(KEYINPUT103), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT103), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n893), .B(new_n912), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n925), .A3(new_n913), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT100), .B1(new_n909), .B2(new_n910), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(new_n921), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n911), .A2(new_n868), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n851), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n893), .B1(new_n928), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n912), .B1(new_n922), .B2(new_n923), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n893), .ZN(new_n935));
  MUX2_X1   g510(.A(new_n932), .B(new_n935), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g511(.A(KEYINPUT104), .B(G1384), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(KEYINPUT68), .A2(KEYINPUT4), .A3(G138), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n471), .B2(new_n472), .ZN(new_n940));
  AOI21_X1  g515(.A(G2105), .B1(new_n940), .B2(new_n490), .ZN(new_n941));
  OAI21_X1  g516(.A(G126), .B1(new_n471), .B2(new_n472), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n462), .B1(new_n942), .B2(new_n495), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n938), .B1(new_n944), .B2(new_n500), .ZN(new_n945));
  INV_X1    g520(.A(new_n475), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(G40), .A3(new_n464), .A4(new_n469), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT46), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n952));
  INV_X1    g527(.A(new_n948), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n709), .B1(KEYINPUT46), .B2(new_n949), .ZN(new_n954));
  INV_X1    g529(.A(G2067), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n754), .B(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT47), .Z(new_n959));
  NAND3_X1  g534(.A1(new_n948), .A2(G1996), .A3(new_n709), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT106), .Z(new_n961));
  OAI21_X1  g536(.A(new_n956), .B1(G1996), .B2(new_n709), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n948), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT107), .ZN(new_n965));
  INV_X1    g540(.A(new_n791), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n785), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n754), .A2(G2067), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n953), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n785), .A2(new_n966), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n948), .B1(new_n971), .B2(new_n967), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n953), .A2(G1986), .A3(G290), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n959), .B(new_n970), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G8), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n501), .A2(KEYINPUT109), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT109), .B1(new_n501), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n470), .A2(new_n982), .A3(new_n475), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n572), .B(G1981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n985), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n989));
  OAI221_X1 g564(.A(new_n984), .B1(new_n985), .B2(new_n986), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n564), .A2(new_n566), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G1981), .B2(new_n572), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(KEYINPUT110), .A3(G1976), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G288), .B2(new_n991), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n984), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n992), .A2(G1976), .ZN(new_n999));
  OR3_X1    g574(.A1(new_n998), .A2(KEYINPUT52), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(KEYINPUT52), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n990), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n501), .A2(new_n978), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n501), .A2(KEYINPUT109), .A3(new_n978), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n947), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2090), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n937), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n983), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n944), .B2(new_n500), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1004), .A2(KEYINPUT108), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(G1971), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n977), .B1(new_n1013), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G166), .A2(new_n977), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT55), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n994), .A2(new_n984), .B1(new_n1003), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT50), .B1(new_n979), .B2(new_n980), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n983), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n699), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1022), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1025), .B1(new_n1032), .B2(G8), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1002), .A2(new_n1033), .A3(new_n1026), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1019), .B1(new_n979), .B2(new_n980), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n983), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1004), .A2(new_n1019), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n983), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n692), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1011), .A2(G2084), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n977), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G168), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT63), .B1(new_n1034), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT63), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n1002), .A2(new_n1045), .A3(new_n1026), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1027), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n555), .A2(new_n1051), .A3(new_n559), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n555), .B2(new_n559), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n947), .B1(new_n945), .B2(KEYINPUT45), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT108), .B1(new_n1004), .B2(new_n1019), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1016), .B(KEYINPUT45), .C1(new_n501), .C2(new_n978), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1056), .B(new_n1057), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1956), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1007), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n743), .B1(new_n1066), .B2(new_n1029), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1060), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(KEYINPUT114), .A3(new_n1055), .ZN(new_n1069));
  INV_X1    g644(.A(G1348), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT50), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1010), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n981), .A2(KEYINPUT113), .A3(new_n955), .A4(new_n983), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1006), .A2(new_n955), .A3(new_n983), .A4(new_n1008), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n591), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1065), .A2(new_n1069), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1067), .A2(new_n1054), .A3(new_n1060), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT117), .B1(new_n1087), .B2(new_n591), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1089), .B(new_n590), .C1(new_n1078), .C2(new_n1086), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1088), .A2(new_n1090), .B1(new_n1086), .B2(new_n1078), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1056), .B(new_n949), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1006), .A2(new_n983), .A3(new_n1008), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n545), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT59), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT114), .B1(new_n1068), .B2(new_n1055), .ZN(new_n1098));
  AOI211_X1 g673(.A(new_n1064), .B(new_n1054), .C1(new_n1067), .C2(new_n1060), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1082), .A2(KEYINPUT61), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1011), .A2(new_n1070), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT60), .B1(new_n1103), .B2(new_n1074), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1089), .B1(new_n1104), .B2(new_n590), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n591), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1068), .B2(new_n1055), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT116), .B(new_n1054), .C1(new_n1067), .C2(new_n1060), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1082), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1091), .A2(new_n1102), .A3(new_n1108), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1085), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(G2078), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n945), .B2(KEYINPUT45), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n1015), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1056), .B(new_n714), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1117), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1011), .B2(new_n680), .ZN(new_n1124));
  AOI211_X1 g699(.A(KEYINPUT120), .B(G1961), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1122), .B(G301), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT121), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n680), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT120), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1011), .A2(new_n1123), .A3(new_n680), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(G301), .A4(new_n1122), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT45), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(new_n947), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(new_n1038), .A3(new_n1036), .A4(new_n1118), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1117), .A2(new_n1121), .B1(new_n1011), .B2(new_n680), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1127), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1145), .A3(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1137), .A2(new_n1138), .A3(G301), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT54), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1122), .B(KEYINPUT123), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1151), .B1(new_n1156), .B2(G171), .ZN(new_n1157));
  AOI211_X1 g732(.A(KEYINPUT124), .B(G301), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT125), .B(new_n1150), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1116), .A2(new_n1147), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n947), .B1(new_n1161), .B2(new_n1019), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1037), .B1(new_n1162), .B2(KEYINPUT112), .ZN(new_n1163));
  AOI21_X1  g738(.A(G1966), .B1(new_n1163), .B2(new_n1136), .ZN(new_n1164));
  OAI211_X1 g739(.A(G8), .B(G286), .C1(new_n1164), .C2(new_n1042), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1044), .A2(KEYINPUT118), .A3(G286), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT51), .B1(new_n1044), .B2(KEYINPUT119), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1136), .A2(new_n1038), .A3(new_n1036), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1042), .B1(new_n1171), .B2(new_n692), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n977), .B1(new_n1172), .B2(G168), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n1172), .B2(new_n977), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1164), .A2(G286), .A3(new_n1042), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1176), .B(KEYINPUT51), .C1(new_n1177), .C2(new_n977), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1169), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT123), .B1(new_n1131), .B2(new_n1122), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1155), .ZN(new_n1181));
  OAI21_X1  g756(.A(G171), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT124), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1156), .A2(new_n1151), .A3(G171), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1149), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1179), .B1(new_n1185), .B2(KEYINPUT125), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1179), .A2(KEYINPUT62), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1169), .A2(new_n1174), .A3(new_n1178), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1140), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1160), .A2(new_n1186), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1050), .B1(new_n1192), .B2(new_n1034), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n948), .A2(G1986), .A3(G290), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n974), .A2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT105), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n973), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n976), .B1(new_n1193), .B2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1200));
  NOR2_X1   g774(.A1(G227), .A2(new_n457), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n637), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1202), .B1(new_n672), .B2(new_n675), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(new_n854), .ZN(new_n1204));
  INV_X1    g778(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1200), .B1(new_n932), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g780(.A(KEYINPUT127), .B(new_n1204), .C1(new_n924), .C2(new_n931), .ZN(new_n1207));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n932), .A2(new_n1205), .ZN(G225));
endmodule


