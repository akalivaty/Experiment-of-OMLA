//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n191), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G137), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT64), .B(new_n203), .C1(new_n199), .C2(G137), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n197), .A2(G134), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT64), .B1(new_n206), .B2(new_n203), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n201), .B(new_n202), .C1(new_n205), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n203), .B1(new_n199), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n202), .B1(new_n213), .B2(new_n201), .ZN(new_n214));
  OAI211_X1 g028(.A(KEYINPUT65), .B(new_n196), .C1(new_n209), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n189), .A3(new_n191), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n193), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n200), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n208), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n201), .B1(new_n205), .B2(new_n207), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n208), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n227), .B2(new_n196), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n187), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR3_X1   g045(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n233));
  INV_X1    g047(.A(G113), .ZN(new_n234));
  OAI22_X1  g048(.A1(new_n231), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n233), .A3(new_n234), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n244), .A2(new_n230), .B1(KEYINPUT2), .B2(G113), .ZN(new_n245));
  INV_X1    g059(.A(new_n240), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n235), .A2(KEYINPUT67), .A3(new_n240), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n196), .B1(new_n209), .B2(new_n214), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(KEYINPUT68), .B(new_n196), .C1(new_n209), .C2(new_n214), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n257), .A2(G128), .B1(new_n189), .B2(new_n191), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n217), .A2(new_n189), .A3(new_n191), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT69), .B(new_n218), .C1(new_n193), .C2(new_n219), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n260), .A2(new_n208), .A3(new_n261), .A4(new_n222), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n254), .A2(KEYINPUT30), .A3(new_n255), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n229), .A2(new_n251), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n254), .A2(new_n250), .A3(new_n255), .A4(new_n262), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT27), .Z(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n255), .A2(new_n262), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT68), .B1(new_n227), .B2(new_n196), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(new_n251), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n208), .A2(new_n220), .A3(new_n222), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n195), .B1(new_n226), .B2(new_n208), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n252), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n250), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT28), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n271), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n251), .A2(new_n277), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT28), .B1(new_n284), .B2(new_n262), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n272), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT71), .B(G902), .Z(new_n290));
  OAI21_X1  g104(.A(new_n251), .B1(new_n273), .B2(new_n274), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n265), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT70), .B(new_n251), .C1(new_n273), .C2(new_n274), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(KEYINPUT29), .A3(new_n283), .A4(new_n286), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n289), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n264), .A2(new_n283), .A3(new_n265), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT31), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n264), .A2(new_n301), .A3(new_n283), .A4(new_n265), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n251), .B1(new_n224), .B2(new_n228), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(new_n265), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n271), .B1(new_n305), .B2(new_n285), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NOR2_X1   g122(.A1(G472), .A2(G902), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n298), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT73), .ZN(new_n317));
  OR3_X1    g131(.A1(new_n315), .A2(KEYINPUT73), .A3(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n190), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n202), .A3(new_n324), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n319), .A2(new_n188), .A3(new_n321), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n202), .B1(new_n332), .B2(new_n324), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT17), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n323), .A2(new_n334), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(KEYINPUT88), .A3(new_n324), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT18), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n202), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n202), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n332), .A2(KEYINPUT88), .A3(new_n342), .A4(new_n324), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n317), .A2(new_n318), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  XNOR2_X1  g160(.A(G125), .B(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n188), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  INV_X1    g165(.A(G104), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n338), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n325), .A2(new_n326), .A3(G131), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(new_n336), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT19), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n317), .B2(new_n318), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n347), .A2(KEYINPUT19), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n188), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n327), .A2(KEYINPUT89), .A3(new_n333), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n357), .A2(new_n323), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT90), .A3(new_n350), .ZN(new_n364));
  INV_X1    g178(.A(new_n353), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT90), .B1(new_n363), .B2(new_n350), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n354), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n369));
  NOR2_X1   g183(.A1(G475), .A2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT91), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n370), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n368), .A2(new_n377), .A3(new_n369), .A4(new_n370), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G902), .ZN(new_n380));
  INV_X1    g194(.A(new_n354), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n353), .B1(new_n338), .B2(new_n350), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G475), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G952), .ZN(new_n386));
  AOI211_X1 g200(.A(G953), .B(new_n386), .C1(G234), .C2(G237), .ZN(new_n387));
  AOI211_X1 g201(.A(new_n330), .B(new_n290), .C1(G234), .C2(G237), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT21), .B(G898), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT15), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G478), .ZN(new_n392));
  INV_X1    g206(.A(G122), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G116), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n238), .A2(G122), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(G128), .A3(new_n190), .ZN(new_n400));
  XNOR2_X1  g214(.A(G128), .B(G143), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n400), .B(G134), .C1(new_n402), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n199), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(KEYINPUT14), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n238), .A3(G122), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT93), .A4(new_n394), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n409), .B(G107), .C1(KEYINPUT93), .C2(new_n408), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n401), .B(new_n199), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n396), .A2(new_n397), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT9), .B(G234), .ZN(new_n414));
  INV_X1    g228(.A(G217), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n414), .A2(new_n415), .A3(G953), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n405), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n405), .B2(new_n413), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n290), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT94), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT94), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n290), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n392), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n419), .A2(KEYINPUT94), .B1(new_n391), .B2(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n385), .A2(new_n390), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(KEYINPUT25), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n216), .A2(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n236), .A2(G128), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT24), .B(G110), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G110), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT23), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n236), .B2(G128), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n431), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT72), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT72), .A4(new_n431), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n434), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n319), .A2(new_n188), .A3(new_n321), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n188), .B1(new_n319), .B2(new_n321), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n432), .A2(new_n433), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n437), .A2(new_n438), .A3(new_n435), .A4(new_n431), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n188), .B2(new_n347), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n323), .A2(KEYINPUT74), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n448), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n348), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n453), .B2(new_n445), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n446), .A2(new_n450), .A3(new_n454), .A4(KEYINPUT75), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n458), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n290), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n429), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n468));
  OAI221_X1 g282(.A(new_n290), .B1(new_n428), .B2(KEYINPUT25), .C1(new_n468), .C2(new_n459), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n415), .B1(new_n290), .B2(G234), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(G902), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n468), .B2(new_n459), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n312), .A2(new_n427), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n220), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n315), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n195), .A2(G125), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(KEYINPUT84), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n330), .A2(G224), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n485), .B(new_n486), .Z(new_n487));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n397), .A3(G104), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT3), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n488), .A2(new_n491), .A3(new_n397), .A4(G104), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n397), .A2(G104), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G101), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n490), .A2(new_n497), .A3(new_n492), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n500), .A3(G101), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n499), .A2(new_n249), .A3(new_n248), .A4(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g317(.A(G113), .B1(new_n237), .B2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n247), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n352), .A2(G107), .ZN(new_n506));
  OAI21_X1  g320(.A(G101), .B1(new_n506), .B2(new_n493), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G110), .B(G122), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(KEYINPUT83), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n509), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT82), .B1(new_n502), .B2(new_n509), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT6), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n487), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n485), .A2(KEYINPUT7), .A3(new_n486), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n508), .B(new_n247), .C1(new_n503), .C2(new_n504), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n510), .B(KEYINPUT8), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(new_n504), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n525), .A2(new_n526), .B1(new_n245), .B2(new_n246), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n522), .B(new_n523), .C1(new_n527), .C2(new_n508), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n481), .A2(new_n482), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n486), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n521), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n380), .B1(new_n532), .B2(new_n512), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n479), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n487), .ZN(new_n535));
  INV_X1    g349(.A(new_n513), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n502), .A2(new_n509), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT82), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n502), .A2(KEYINPUT82), .A3(new_n509), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n511), .B1(new_n541), .B2(KEYINPUT6), .ZN(new_n542));
  INV_X1    g356(.A(new_n519), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n533), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n478), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n534), .A2(new_n546), .A3(KEYINPUT86), .ZN(new_n547));
  OAI21_X1  g361(.A(G214), .B1(G237), .B2(G902), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n544), .A2(new_n549), .A3(new_n545), .A4(new_n478), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n260), .A2(new_n261), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n498), .A2(KEYINPUT10), .A3(new_n507), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n498), .A2(KEYINPUT10), .A3(new_n507), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(KEYINPUT80), .A3(new_n260), .A4(new_n261), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n227), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n257), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n189), .A2(KEYINPUT79), .A3(KEYINPUT1), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(G128), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n193), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n259), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n561), .B1(new_n567), .B2(new_n508), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n499), .A2(new_n501), .A3(new_n196), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n559), .A2(new_n560), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G140), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n330), .A2(G227), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n567), .A2(new_n508), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n220), .B1(new_n498), .B2(new_n507), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT81), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n227), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT12), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n480), .A2(new_n508), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n508), .B2(new_n567), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n578), .A3(new_n583), .A4(new_n227), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n570), .A2(new_n574), .A3(new_n580), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n556), .A2(new_n558), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n569), .A2(new_n568), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n227), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n574), .B1(new_n589), .B2(new_n570), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n552), .B(new_n290), .C1(new_n586), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(G469), .A2(G902), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n587), .A2(new_n227), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n580), .A2(new_n584), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n573), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n589), .A2(new_n570), .A3(new_n574), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(G469), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G221), .B1(new_n414), .B2(G902), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT77), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n551), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n477), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n307), .A2(new_n309), .ZN(new_n606));
  INV_X1    g420(.A(G472), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n307), .B2(new_n290), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n608), .B2(KEYINPUT95), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n610), .B(new_n607), .C1(new_n307), .C2(new_n290), .ZN(new_n611));
  NOR4_X1   g425(.A1(new_n609), .A2(new_n611), .A3(new_n475), .A4(new_n602), .ZN(new_n612));
  INV_X1    g426(.A(new_n548), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n534), .B2(new_n546), .ZN(new_n614));
  INV_X1    g428(.A(new_n390), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n417), .A2(new_n418), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(KEYINPUT96), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(KEYINPUT96), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI22_X1  g434(.A1(new_n417), .A2(new_n418), .B1(KEYINPUT96), .B2(new_n617), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(G478), .A3(new_n290), .A4(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n419), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n379), .B2(new_n384), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n614), .A2(new_n615), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n612), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  OAI21_X1  g446(.A(KEYINPUT99), .B1(new_n373), .B2(new_n375), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n368), .A2(new_n634), .A3(new_n370), .A4(new_n374), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT98), .B1(new_n373), .B2(new_n375), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  AOI211_X1 g451(.A(new_n637), .B(new_n374), .C1(new_n368), .C2(new_n370), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n633), .B(new_n635), .C1(new_n636), .C2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n384), .A2(KEYINPUT100), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n383), .B2(G475), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n425), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n615), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  INV_X1    g461(.A(new_n614), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n612), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n464), .A2(KEYINPUT36), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n463), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n463), .A2(new_n653), .ZN(new_n655));
  INV_X1    g469(.A(new_n473), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n470), .B2(new_n471), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n385), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n615), .A4(new_n425), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n661), .A2(new_n609), .A3(new_n611), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n603), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n387), .B1(new_n388), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n639), .A2(new_n643), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n602), .A2(new_n658), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n312), .A2(new_n614), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NAND2_X1  g486(.A1(new_n547), .A2(new_n550), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT38), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT38), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n547), .A2(new_n675), .A3(new_n550), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n425), .B1(new_n379), .B2(new_n384), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n548), .A3(new_n658), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n293), .A2(new_n294), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n680), .B2(new_n271), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n266), .A2(new_n283), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n607), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n310), .B2(new_n311), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n667), .B(KEYINPUT39), .Z(new_n686));
  NAND3_X1  g500(.A1(new_n598), .A2(new_n601), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n598), .A2(new_n689), .A3(new_n601), .A4(new_n686), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n679), .A2(new_n685), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT102), .B1(new_n677), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n548), .A3(new_n658), .A4(new_n678), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n606), .A2(KEYINPUT32), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n683), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n570), .A2(new_n574), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n570), .A2(new_n580), .A3(new_n584), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n697), .A2(new_n589), .B1(new_n698), .B2(new_n573), .ZN(new_n699));
  OAI21_X1  g513(.A(G469), .B1(new_n699), .B2(G902), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n600), .B1(new_n700), .B2(new_n591), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n689), .B1(new_n701), .B2(new_n686), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n693), .A2(new_n696), .A3(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n547), .A2(new_n675), .A3(new_n550), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n675), .B1(new_n547), .B2(new_n550), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n692), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n190), .ZN(G45));
  AOI211_X1 g524(.A(new_n667), .B(new_n626), .C1(new_n379), .C2(new_n384), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n312), .A2(new_n614), .A3(new_n670), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  INV_X1    g527(.A(new_n599), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n290), .B1(new_n586), .B2(new_n590), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n591), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(KEYINPUT103), .A3(G469), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n312), .A2(new_n476), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n628), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND2_X1  g538(.A1(new_n649), .A2(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND2_X1  g540(.A1(new_n694), .A2(new_n695), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n661), .B1(new_n727), .B2(new_n298), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n720), .A2(new_n614), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n295), .A2(new_n286), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n732), .B(new_n300), .C1(new_n733), .C2(new_n283), .ZN(new_n734));
  INV_X1    g548(.A(new_n300), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n283), .B1(new_n295), .B2(new_n286), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT104), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n737), .A3(new_n302), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n608), .B(new_n475), .C1(new_n309), .C2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n614), .A2(new_n615), .A3(new_n678), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n741), .A3(KEYINPUT105), .A4(new_n720), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n309), .ZN(new_n744));
  INV_X1    g558(.A(new_n608), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n720), .A3(new_n476), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n743), .B1(new_n746), .B2(new_n740), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NAND3_X1  g563(.A1(new_n744), .A2(new_n745), .A3(new_n659), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n720), .A2(new_n614), .A3(new_n711), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n315), .ZN(G27));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n613), .B1(new_n547), .B2(new_n550), .ZN(new_n755));
  INV_X1    g569(.A(new_n588), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n560), .B1(new_n756), .B2(new_n559), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n573), .B1(new_n593), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g572(.A(G469), .B(new_n466), .C1(new_n758), .C2(new_n585), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n597), .A2(new_n592), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n599), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n312), .A3(new_n476), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n711), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n754), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n613), .B(new_n761), .C1(new_n547), .C2(new_n550), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n475), .B1(new_n727), .B2(new_n298), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT42), .A4(new_n711), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n767), .A3(new_n669), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n385), .B2(new_n626), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n385), .B(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n625), .A2(KEYINPUT43), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n659), .B1(new_n609), .B2(new_n611), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT44), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n777), .A2(new_n779), .A3(new_n782), .A4(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n595), .A2(new_n596), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n595), .A2(KEYINPUT45), .A3(new_n596), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(G469), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n592), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n759), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT106), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(new_n793), .A3(KEYINPUT46), .A4(new_n592), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n592), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT106), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n599), .A2(new_n797), .A3(new_n686), .A4(new_n755), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  INV_X1    g613(.A(new_n774), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n385), .B(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n776), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n799), .B1(new_n804), .B2(new_n778), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n784), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT109), .B(G137), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G39));
  INV_X1    g623(.A(new_n755), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n810), .A2(new_n312), .A3(new_n764), .A4(new_n476), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n599), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT47), .B1(new_n797), .B2(new_n599), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  NAND2_X1  g629(.A1(new_n777), .A2(new_n387), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT115), .Z(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n810), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n721), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT48), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n817), .A2(new_n648), .A3(new_n746), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT117), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n476), .A2(new_n387), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n696), .A3(new_n720), .A4(new_n755), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n386), .B(G953), .C1(new_n825), .C2(new_n627), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n820), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n608), .B(new_n658), .C1(new_n738), .C2(new_n309), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n818), .A2(new_n720), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n825), .A2(new_n660), .A3(new_n626), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT116), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n812), .A2(new_n813), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n718), .A2(new_n719), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n601), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n818), .B(new_n739), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n817), .ZN(new_n839));
  INV_X1    g653(.A(new_n746), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n613), .A3(new_n677), .A4(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT50), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n828), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n841), .B(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n833), .A3(KEYINPUT51), .A4(new_n837), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n827), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n385), .A2(new_n425), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n615), .B1(new_n848), .B2(new_n627), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n551), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n649), .A2(new_n721), .B1(new_n850), .B2(new_n612), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n728), .A2(new_n729), .B1(new_n477), .B2(new_n603), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n662), .A2(new_n603), .B1(new_n721), .B2(new_n628), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n748), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n829), .A2(new_n766), .A3(new_n711), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n426), .A2(new_n642), .A3(new_n640), .A4(new_n667), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(new_n639), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n755), .A2(new_n857), .A3(new_n312), .A4(new_n670), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n855), .A2(new_n771), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(new_n769), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n854), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n748), .A2(new_n852), .A3(new_n851), .A4(new_n853), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n769), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT110), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n671), .B1(new_n750), .B2(new_n751), .ZN(new_n867));
  INV_X1    g681(.A(new_n657), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n667), .B(KEYINPUT113), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n472), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n761), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n685), .A3(new_n614), .A4(new_n678), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n712), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n867), .A2(new_n873), .A3(KEYINPUT52), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT52), .B1(new_n867), .B2(new_n873), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n671), .B(KEYINPUT112), .C1(new_n750), .C2(new_n751), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n712), .A3(new_n872), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT52), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n879), .B1(new_n884), .B2(new_n875), .ZN(new_n885));
  AOI211_X1 g699(.A(KEYINPUT114), .B(new_n874), .C1(new_n883), .C2(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n854), .A2(new_n860), .A3(KEYINPUT53), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n878), .A2(new_n888), .A3(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n861), .B1(new_n854), .B2(new_n860), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT110), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT111), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n885), .A2(new_n886), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT111), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n862), .A2(new_n895), .A3(new_n865), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n866), .A2(new_n877), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT53), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(KEYINPUT54), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n889), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n847), .A2(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n835), .B(KEYINPUT49), .Z(new_n903));
  NAND4_X1  g717(.A1(new_n476), .A2(new_n548), .A3(new_n601), .A4(new_n625), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n904), .A2(new_n775), .A3(new_n685), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n677), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n906), .ZN(G75));
  OAI211_X1 g721(.A(new_n479), .B(new_n466), .C1(new_n878), .C2(new_n888), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n542), .A2(new_n543), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT118), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n535), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n908), .A2(new_n909), .A3(new_n914), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n330), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT119), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n916), .A2(new_n922), .A3(new_n917), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(G51));
  OAI21_X1  g738(.A(KEYINPUT54), .B1(new_n878), .B2(new_n888), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n889), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n592), .B(KEYINPUT57), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n590), .B2(new_n586), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n878), .A2(new_n888), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n466), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n931), .A2(new_n789), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n918), .B1(new_n929), .B2(new_n932), .ZN(G54));
  INV_X1    g747(.A(new_n368), .ZN(new_n934));
  NAND2_X1  g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n919), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G60));
  NAND2_X1  g753(.A1(new_n620), .A2(new_n621), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n926), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n901), .B2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n918), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT60), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n930), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n465), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n654), .A2(new_n655), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n930), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n919), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n950), .A2(new_n919), .A3(new_n952), .A4(new_n954), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(new_n389), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n330), .B1(new_n959), .B2(G224), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n863), .B2(new_n330), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n912), .B1(G898), .B2(new_n330), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n961), .B(new_n962), .Z(G69));
  AOI21_X1  g777(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n767), .A2(new_n614), .A3(new_n678), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(new_n599), .A3(new_n686), .A4(new_n797), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n814), .A2(new_n966), .A3(new_n769), .A4(new_n771), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n798), .A2(new_n805), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n783), .B2(new_n781), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n881), .A2(new_n712), .A3(new_n882), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT123), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  INV_X1    g786(.A(new_n712), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n867), .B2(new_n880), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n807), .A2(new_n972), .A3(new_n882), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n967), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n330), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n229), .A2(new_n263), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT121), .Z(new_n979));
  OR2_X1    g793(.A1(new_n359), .A2(new_n360), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(new_n981));
  OAI211_X1 g795(.A(new_n977), .B(new_n981), .C1(new_n666), .C2(new_n330), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n964), .B1(new_n982), .B2(KEYINPUT122), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n970), .B2(new_n709), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n692), .A2(new_n708), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(KEYINPUT62), .A3(new_n882), .A4(new_n974), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n767), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n848), .A2(new_n627), .ZN(new_n990));
  OR4_X1    g804(.A1(new_n989), .A2(new_n810), .A3(new_n687), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n814), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n784), .B2(new_n806), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n982), .B1(new_n995), .B2(new_n981), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n983), .B(new_n996), .Z(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n976), .B2(new_n854), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n266), .A2(new_n283), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n919), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n988), .A2(new_n854), .A3(new_n993), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(KEYINPUT124), .A3(new_n999), .ZN(new_n1006));
  INV_X1    g820(.A(new_n682), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(KEYINPUT124), .B1(new_n1005), .B2(new_n999), .ZN(new_n1009));
  OAI21_X1  g823(.A(KEYINPUT125), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1005), .A2(new_n999), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT125), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n1014), .A3(new_n1007), .A4(new_n1006), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1004), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1007), .A2(new_n1002), .A3(new_n1000), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n897), .A2(new_n899), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n897), .A2(new_n1020), .A3(new_n899), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1016), .A2(new_n1022), .A3(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(G57));
endmodule


