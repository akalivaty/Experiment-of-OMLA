//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968;
  OR3_X1    g000(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n202), .A2(KEYINPUT94), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT94), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n202), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n205), .A3(new_n208), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n210), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT95), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT17), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(KEYINPUT16), .A3(new_n227), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G8gat), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n232), .A3(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(KEYINPUT96), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT96), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n237), .A3(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n219), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n219), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n243), .A3(new_n238), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n241), .B(KEYINPUT13), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n225), .A2(new_n234), .B1(new_n219), .B2(new_n239), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n241), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT11), .ZN(new_n255));
  INV_X1    g054(.A(G169gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n248), .B(new_n253), .C1(KEYINPUT98), .C2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT99), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n242), .A2(KEYINPUT98), .A3(new_n247), .ZN(new_n263));
  INV_X1    g062(.A(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n247), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n252), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n262), .B1(new_n261), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT34), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n274));
  INV_X1    g073(.A(G113gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(G120gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(G120gat), .ZN(new_n277));
  INV_X1    g076(.A(G120gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(G113gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n287), .B2(new_n277), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290));
  INV_X1    g089(.A(G134gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G127gat), .ZN(new_n292));
  INV_X1    g091(.A(G127gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G134gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT70), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT71), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n291), .A2(G127gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT70), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n290), .B1(new_n293), .B2(G134gat), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n289), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n306));
  OAI211_X1 g105(.A(KEYINPUT71), .B(new_n297), .C1(new_n284), .C2(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n289), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n286), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n319));
  AND4_X1   g118(.A1(KEYINPUT25), .A2(new_n313), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT24), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(G183gat), .A3(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT67), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n325), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n320), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n312), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n313), .A3(new_n318), .A4(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n326), .A2(KEYINPUT64), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n326), .A2(KEYINPUT64), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n338), .A2(new_n339), .B1(new_n322), .B2(new_n324), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n333), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  INV_X1    g142(.A(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(KEYINPUT28), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n345), .B(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n316), .A2(new_n317), .B1(new_n352), .B2(new_n312), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n351), .A2(new_n353), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n311), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n309), .B1(new_n308), .B2(new_n289), .ZN(new_n358));
  AOI211_X1 g157(.A(KEYINPUT72), .B(new_n288), .C1(new_n306), .C2(new_n307), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n285), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n332), .A2(new_n341), .B1(new_n348), .B2(new_n354), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n273), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT76), .B(new_n273), .C1(new_n357), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT34), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT75), .B1(new_n357), .B2(new_n362), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n311), .A2(new_n356), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n360), .A2(new_n361), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n272), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n367), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n272), .A3(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(KEYINPUT32), .ZN(new_n379));
  XOR2_X1   g178(.A(G15gat), .B(G43gat), .Z(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n382), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n376), .B(KEYINPUT32), .C1(new_n377), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT77), .B1(new_n375), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n371), .B1(new_n370), .B2(new_n372), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n271), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(KEYINPUT34), .B1(new_n365), .B2(new_n366), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n385), .A4(new_n383), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(KEYINPUT34), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n367), .B1(new_n385), .B2(new_n383), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT36), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT36), .ZN(new_n399));
  AOI211_X1 g198(.A(new_n399), .B(new_n396), .C1(new_n387), .C2(new_n393), .ZN(new_n400));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n342), .B2(new_n355), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(KEYINPUT79), .B(KEYINPUT29), .Z(new_n404));
  OAI21_X1  g203(.A(new_n401), .B1(new_n361), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(G211gat), .A2(G218gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(G211gat), .A2(G218gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  INV_X1    g210(.A(G197gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(G204gat), .ZN(new_n413));
  INV_X1    g212(.A(G204gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(G197gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(G197gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(G204gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n407), .A2(KEYINPUT22), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n410), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n409), .B(new_n421), .C1(new_n416), .C2(new_n419), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n401), .B1(new_n361), .B2(KEYINPUT29), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT78), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT78), .B1(new_n417), .B2(new_n418), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n409), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n420), .A2(new_n410), .A3(new_n422), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n403), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT30), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n439), .A2(KEYINPUT30), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n434), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n437), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G141gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(G148gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT80), .B(G141gat), .ZN(new_n453));
  INV_X1    g252(.A(G148gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT2), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G155gat), .ZN(new_n459));
  INV_X1    g258(.A(G162gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n454), .A2(G141gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n457), .B1(new_n451), .B2(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G155gat), .B(G162gat), .Z(new_n464));
  AOI22_X1  g263(.A1(new_n455), .A2(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n360), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n465), .B(new_n285), .C1(new_n358), .C2(new_n359), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G225gat), .A2(G233gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n465), .B(KEYINPUT3), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n360), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT4), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n311), .B2(new_n465), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT81), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n311), .A2(new_n476), .A3(new_n465), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n475), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n473), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n311), .A2(new_n487), .A3(new_n476), .A4(new_n465), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT82), .B1(new_n468), .B2(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n478), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n360), .A2(new_n474), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n470), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n449), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n469), .B2(new_n471), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n483), .A2(new_n484), .A3(new_n475), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n484), .B1(new_n483), .B2(new_n475), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n448), .A3(new_n493), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT6), .B(new_n449), .C1(new_n486), .C2(new_n494), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n444), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n423), .B2(new_n424), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n465), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n404), .B1(new_n465), .B2(new_n507), .ZN(new_n509));
  OAI211_X1 g308(.A(G228gat), .B(G233gat), .C1(new_n509), .C2(new_n433), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT85), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G228gat), .A2(G233gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n455), .A2(new_n461), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n463), .A2(new_n464), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n404), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n517), .B2(new_n425), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT3), .B1(new_n433), .B2(new_n505), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n518), .B(new_n519), .C1(new_n465), .C2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n516), .B1(new_n423), .B2(new_n424), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n465), .B1(new_n522), .B2(new_n507), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n509), .A2(new_n433), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n512), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n511), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G22gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  INV_X1    g327(.A(G22gat), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n511), .A2(new_n521), .A3(new_n525), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532));
  XNOR2_X1  g331(.A(G78gat), .B(G106gat), .ZN(new_n533));
  INV_X1    g332(.A(G50gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT84), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n532), .B1(new_n531), .B2(new_n538), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n527), .A2(new_n530), .ZN(new_n541));
  OAI22_X1  g340(.A1(new_n539), .A2(new_n540), .B1(new_n528), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n538), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT87), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n541), .A2(new_n528), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n398), .A2(new_n400), .B1(new_n504), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT40), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n470), .B1(new_n490), .B2(new_n492), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT88), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n467), .A2(new_n556), .A3(new_n468), .A4(new_n470), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT39), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n448), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT39), .B(new_n470), .C1(new_n490), .C2(new_n492), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n561), .A2(new_n495), .A3(new_n444), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n559), .A2(new_n552), .A3(new_n560), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n562), .A2(new_n563), .B1(new_n547), .B2(new_n542), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n503), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n499), .A2(new_n493), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n567), .A2(KEYINPUT91), .A3(KEYINPUT6), .A4(new_n449), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n356), .A2(new_n516), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n402), .B1(new_n571), .B2(new_n401), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n434), .B(new_n570), .C1(new_n572), .C2(new_n433), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n573), .A2(new_n437), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n442), .A2(KEYINPUT37), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n403), .A2(new_n427), .A3(new_n425), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(KEYINPUT37), .C1(new_n572), .C2(new_n425), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n573), .A2(new_n578), .A3(new_n437), .A4(new_n569), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n439), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n502), .A2(new_n566), .A3(new_n568), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n551), .B1(new_n564), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n563), .A2(new_n495), .A3(new_n444), .A4(new_n561), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n582), .A2(new_n548), .A3(new_n584), .A4(new_n551), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n550), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n396), .B1(new_n387), .B2(new_n393), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n444), .A2(KEYINPUT35), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n548), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n502), .A2(new_n566), .A3(new_n568), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n504), .A2(new_n548), .A3(new_n588), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(KEYINPUT35), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n270), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  XOR2_X1   g395(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n597));
  INV_X1    g396(.A(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(G57gat), .ZN(new_n599));
  INV_X1    g398(.A(G57gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT9), .ZN(new_n603));
  AND2_X1   g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT100), .B1(new_n600), .B2(G64gat), .ZN(new_n608));
  MUX2_X1   g407(.A(KEYINPUT100), .B(new_n608), .S(new_n599), .Z(new_n609));
  AOI21_X1  g408(.A(new_n604), .B1(KEYINPUT9), .B2(new_n605), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n615), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n597), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n239), .B1(KEYINPUT21), .B2(new_n612), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n613), .B(new_n614), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n616), .ZN(new_n625));
  INV_X1    g424(.A(new_n597), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n618), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n623), .B1(new_n621), .B2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n596), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n627), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n626), .B1(new_n625), .B2(new_n618), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n622), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n596), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(G85gat), .ZN(new_n640));
  INV_X1    g439(.A(G92gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT7), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n640), .B2(new_n641), .ZN(new_n644));
  NAND3_X1  g443(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G99gat), .B(G106gat), .Z(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n225), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  AND2_X1   g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n652), .A2(new_n219), .B1(KEYINPUT41), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n651), .B2(new_n654), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n638), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(G134gat), .B(G162gat), .Z(new_n660));
  NOR2_X1   g459(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n659), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n637), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n612), .A2(new_n650), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT102), .B1(new_n646), .B2(new_n647), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n649), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n647), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n611), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n652), .A2(new_n612), .A3(KEYINPUT10), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n666), .A2(new_n670), .A3(new_n674), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G120gat), .B(G148gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n673), .A2(KEYINPUT104), .A3(new_n674), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n676), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n683), .B1(new_n687), .B2(new_n682), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT105), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n690), .B(new_n683), .C1(new_n687), .C2(new_n682), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n664), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n595), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n502), .A2(new_n503), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n227), .ZN(G1324gat));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND4_X1  g497(.A1(new_n595), .A2(new_n444), .A3(new_n693), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(KEYINPUT42), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(KEYINPUT42), .ZN(new_n702));
  INV_X1    g501(.A(new_n444), .ZN(new_n703));
  OAI21_X1  g502(.A(G8gat), .B1(new_n694), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT107), .ZN(G1325gat));
  NOR2_X1   g505(.A1(new_n398), .A2(new_n400), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n694), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n588), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(G15gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n694), .B2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n694), .A2(new_n548), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT108), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n714), .B(new_n715), .Z(G1327gat));
  INV_X1    g515(.A(new_n637), .ZN(new_n717));
  INV_X1    g516(.A(new_n663), .ZN(new_n718));
  INV_X1    g517(.A(new_n692), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n595), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G29gat), .A3(new_n695), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT45), .Z(new_n722));
  NAND3_X1  g521(.A1(new_n582), .A2(new_n548), .A3(new_n584), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT92), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n549), .B1(new_n724), .B2(new_n585), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n718), .C1(new_n725), .C2(new_n593), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n261), .A2(new_n266), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n637), .A2(new_n692), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n593), .B1(new_n725), .B2(KEYINPUT109), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n587), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n663), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n726), .B(new_n729), .C1(new_n733), .C2(KEYINPUT44), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n695), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n722), .A2(new_n735), .ZN(G1328gat));
  NOR3_X1   g535(.A1(new_n720), .A2(G36gat), .A3(new_n703), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n734), .B2(new_n703), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  NAND2_X1  g539(.A1(new_n707), .A2(G43gat), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n720), .A2(new_n710), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n734), .A2(new_n741), .B1(new_n742), .B2(G43gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1330gat));
  OAI21_X1  g544(.A(new_n534), .B1(new_n720), .B2(new_n548), .ZN(new_n746));
  INV_X1    g545(.A(new_n548), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n734), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n732), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n637), .A2(new_n728), .A3(new_n663), .A4(new_n692), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n695), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n444), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n759), .B2(new_n758), .ZN(G1333gat));
  NAND2_X1  g561(.A1(new_n754), .A2(new_n588), .ZN(new_n763));
  INV_X1    g562(.A(G71gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n708), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n763), .A2(new_n764), .B1(new_n754), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n754), .A2(new_n747), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g569(.A1(new_n717), .A2(new_n728), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n719), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n726), .B(new_n772), .C1(new_n733), .C2(KEYINPUT44), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n773), .A2(new_n640), .A3(new_n695), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n771), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n751), .A2(new_n718), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n779), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n733), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n780), .A2(new_n755), .A3(new_n692), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n774), .B1(new_n640), .B2(new_n783), .ZN(G1336gat));
  NOR2_X1   g583(.A1(new_n703), .A2(G92gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n780), .A2(new_n692), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n773), .B2(new_n703), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT52), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n786), .B(new_n787), .C1(KEYINPUT113), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n773), .B2(new_n708), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n710), .A2(new_n719), .A3(G99gat), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n782), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(G1338gat));
  NOR2_X1   g597(.A1(new_n548), .A2(G106gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n692), .A3(new_n782), .A4(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G106gat), .B1(new_n773), .B2(new_n548), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n800), .B(new_n801), .C1(new_n803), .C2(KEYINPUT53), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(new_n683), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n673), .B2(new_n674), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n671), .A2(G230gat), .A3(G233gat), .A4(new_n672), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n682), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n685), .A2(new_n686), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n813), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n809), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT55), .B(new_n813), .C1(new_n814), .C2(new_n816), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n727), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n248), .A2(new_n253), .A3(new_n260), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n251), .A2(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n258), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT117), .B1(new_n823), .B2(new_n258), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n691), .B2(new_n689), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n663), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n819), .A2(new_n820), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n663), .A3(new_n826), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n637), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n664), .A2(new_n727), .A3(new_n692), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT118), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n693), .A2(new_n728), .ZN(new_n835));
  INV_X1    g634(.A(new_n826), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n692), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n727), .A2(new_n819), .A3(new_n820), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n718), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n717), .B1(new_n839), .B2(new_n830), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n695), .A2(new_n444), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n747), .A2(new_n710), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n275), .B1(new_n847), .B2(new_n728), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n269), .A2(G113gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT119), .ZN(G1340gat));
  NOR2_X1   g650(.A1(new_n847), .A2(new_n719), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n278), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n847), .A2(new_n717), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(new_n293), .ZN(G1342gat));
  AOI21_X1  g654(.A(new_n663), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n845), .A2(new_n846), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n857), .B(new_n858), .Z(G1343gat));
  NOR2_X1   g658(.A1(new_n707), .A2(new_n548), .ZN(new_n860));
  AND4_X1   g659(.A1(new_n450), .A2(new_n845), .A3(new_n269), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n862));
  INV_X1    g661(.A(new_n453), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n819), .A2(new_n864), .A3(new_n820), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n819), .B2(new_n820), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n269), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n718), .B1(new_n867), .B2(new_n837), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n717), .B1(new_n868), .B2(new_n830), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT122), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n717), .C1(new_n868), .C2(new_n830), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n835), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n548), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n834), .A2(new_n842), .A3(new_n747), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n873), .A2(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n708), .A2(new_n844), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n878), .A2(new_n270), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n862), .B1(new_n863), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n872), .A2(new_n835), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n829), .A2(KEYINPUT121), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n819), .A2(new_n864), .A3(new_n820), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n827), .B1(new_n887), .B2(new_n269), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n831), .B1(new_n888), .B2(new_n718), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n871), .B1(new_n889), .B2(new_n717), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n875), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n877), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n879), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT123), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n883), .A2(new_n894), .A3(new_n727), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n861), .B1(new_n895), .B2(new_n453), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n881), .B1(new_n896), .B2(new_n897), .ZN(G1344gat));
  NOR3_X1   g697(.A1(new_n719), .A2(G148gat), .A3(new_n444), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n843), .A2(new_n755), .A3(new_n860), .A4(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G148gat), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n893), .A2(KEYINPUT123), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n882), .B(new_n879), .C1(new_n891), .C2(new_n892), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n905), .B2(new_n692), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n889), .A2(new_n717), .B1(new_n270), .B2(new_n693), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n874), .B1(new_n907), .B2(new_n548), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n876), .B2(new_n877), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n909), .A2(new_n708), .A3(new_n692), .A4(new_n844), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n901), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n900), .B1(new_n906), .B2(new_n911), .ZN(G1345gat));
  AND2_X1   g711(.A1(new_n845), .A2(new_n860), .ZN(new_n913));
  AOI21_X1  g712(.A(G155gat), .B1(new_n913), .B2(new_n637), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n637), .A2(G155gat), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT124), .Z(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n905), .B2(new_n916), .ZN(G1346gat));
  NAND3_X1  g716(.A1(new_n913), .A2(new_n460), .A3(new_n718), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n903), .A2(new_n904), .A3(new_n663), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n460), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n755), .A2(new_n703), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n843), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(new_n846), .ZN(new_n923));
  AOI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n727), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n846), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n256), .A3(new_n270), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n924), .A2(new_n926), .ZN(G1348gat));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n692), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(G176gat), .ZN(G1349gat));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n923), .A2(new_n343), .A3(new_n637), .ZN(new_n931));
  OAI21_X1  g730(.A(G183gat), .B1(new_n925), .B2(new_n717), .ZN(new_n932));
  AOI211_X1 g731(.A(new_n930), .B(KEYINPUT60), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n935));
  AND4_X1   g734(.A1(new_n931), .A2(new_n932), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n933), .A2(new_n936), .ZN(G1350gat));
  NAND2_X1  g736(.A1(new_n923), .A2(new_n718), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(G190gat), .ZN(new_n941));
  OAI21_X1  g740(.A(G190gat), .B1(new_n925), .B2(new_n663), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n942), .B2(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n923), .A2(new_n344), .A3(new_n718), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  AND2_X1   g746(.A1(new_n922), .A2(new_n860), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948), .B2(new_n727), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n708), .A2(new_n921), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT127), .Z(new_n951));
  AND2_X1   g750(.A1(new_n909), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n270), .A2(new_n412), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  AND4_X1   g753(.A1(new_n414), .A2(new_n922), .A3(new_n692), .A4(new_n860), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n952), .A2(new_n692), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n414), .ZN(G1353gat));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n708), .A2(new_n637), .A3(new_n921), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n959), .B1(new_n909), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT63), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n959), .A3(new_n637), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1354gat));
  INV_X1    g764(.A(G218gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n966), .A3(new_n718), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n952), .A2(new_n718), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n966), .ZN(G1355gat));
endmodule


