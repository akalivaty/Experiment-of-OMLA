//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT68), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G221), .A3(G220), .A4(G218), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(new_n471), .B2(new_n472), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(G136), .B2(new_n473), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n473), .A2(new_n486), .A3(G138), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n478), .C1(new_n462), .C2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(G126), .B2(new_n479), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(G50), .A2(G543), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g074(.A(G543), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G543), .C1(new_n498), .C2(new_n499), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XOR2_X1   g082(.A(KEYINPUT74), .B(G88), .Z(new_n508));
  OAI21_X1  g083(.A(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(KEYINPUT70), .B(new_n510), .C1(new_n511), .C2(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT6), .B1(new_n511), .B2(KEYINPUT70), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n507), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n521), .A2(new_n522), .A3(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n522), .B1(new_n521), .B2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(new_n502), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n503), .B1(new_n534), .B2(new_n505), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(new_n517), .A3(new_n501), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n540), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n539), .A2(G51), .A3(G543), .A4(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n535), .A2(G63), .A3(G651), .A4(new_n501), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(KEYINPUT77), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n538), .B1(new_n545), .B2(new_n547), .ZN(G168));
  NAND4_X1  g123(.A1(new_n539), .A2(G52), .A3(G543), .A4(new_n541), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n535), .A2(G90), .A3(new_n517), .A4(new_n501), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n501), .A2(G64), .A3(new_n504), .A4(new_n506), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n511), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n507), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n539), .A2(G543), .A3(new_n541), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n561), .A2(new_n562), .B1(new_n536), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT78), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n539), .A2(G53), .A3(G543), .A4(new_n541), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n507), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n517), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n507), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n576), .A2(G651), .B1(new_n578), .B2(G91), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n573), .A2(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n552), .A2(new_n553), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n582), .A2(new_n583), .A3(new_n549), .A4(new_n550), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT79), .B1(new_n551), .B2(new_n554), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G301));
  INV_X1    g162(.A(new_n538), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n546), .B1(new_n542), .B2(new_n543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G286));
  AND3_X1   g166(.A1(new_n539), .A2(G543), .A3(new_n541), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G49), .ZN(new_n593));
  INV_X1    g168(.A(new_n507), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n594), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n578), .A2(G87), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND3_X1  g172(.A1(new_n535), .A2(G61), .A3(new_n501), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n501), .A2(G86), .A3(new_n504), .A4(new_n506), .ZN(new_n602));
  NAND2_X1  g177(.A1(G48), .A2(G543), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n577), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n594), .A2(G60), .ZN(new_n607));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n511), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT80), .B(G47), .Z(new_n610));
  INV_X1    g185(.A(G85), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n561), .A2(new_n610), .B1(new_n536), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND3_X1  g189(.A1(new_n578), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n536), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n507), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(G651), .A2(new_n622), .B1(new_n592), .B2(G54), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n586), .ZN(G284));
  AOI21_X1  g201(.A(new_n625), .B1(G868), .B2(new_n586), .ZN(G321));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI21_X1  g203(.A(KEYINPUT81), .B1(new_n628), .B2(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  MUX2_X1   g205(.A(KEYINPUT81), .B(new_n629), .S(new_n630), .Z(G297));
  MUX2_X1   g206(.A(KEYINPUT81), .B(new_n629), .S(new_n630), .Z(G280));
  INV_X1    g207(.A(new_n624), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G559), .Z(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(G860), .B2(new_n634), .ZN(G148));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n473), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n479), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n478), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT84), .B(G2100), .Z(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n651), .A3(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT85), .Z(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n658), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT90), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n685), .A2(new_n688), .A3(new_n692), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  XNOR2_X1  g277(.A(KEYINPUT30), .B(G28), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OR2_X1    g279(.A1(KEYINPUT31), .A2(G11), .ZN(new_n705));
  NAND2_X1  g280(.A1(KEYINPUT31), .A2(G11), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n644), .B2(new_n704), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT25), .ZN(new_n710));
  INV_X1    g285(.A(new_n464), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n711), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n478), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n710), .B(new_n713), .C1(G139), .C2(new_n473), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(new_n704), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n704), .B2(G33), .ZN(new_n716));
  INV_X1    g291(.A(G2072), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n708), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n473), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n479), .A2(G129), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G32), .B(new_n724), .S(G29), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT27), .B(G1996), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n718), .B1(new_n719), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n704), .B1(new_n729), .B2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(G34), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G160), .B2(G29), .ZN(new_n732));
  AOI22_X1  g307(.A1(G2084), .A2(new_n732), .B1(new_n725), .B2(new_n726), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n733), .B1(G2084), .B2(new_n732), .C1(new_n716), .C2(new_n717), .ZN(new_n734));
  NOR2_X1   g309(.A1(G164), .A2(new_n704), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G27), .B2(new_n704), .ZN(new_n736));
  INV_X1    g311(.A(G2078), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n727), .A2(new_n719), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR4_X1   g316(.A1(new_n728), .A2(new_n734), .A3(new_n738), .A4(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G35), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G162), .B2(G29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT29), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n742), .B1(G1961), .B2(new_n745), .C1(G2090), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G168), .A2(G16), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT96), .B2(new_n750), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1966), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n745), .A2(G1961), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT97), .Z(new_n755));
  NOR3_X1   g330(.A1(new_n749), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n743), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n633), .B2(new_n743), .ZN(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n704), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  OAI21_X1  g337(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n763));
  INV_X1    g338(.A(G116), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  AOI22_X1  g341(.A1(G128), .A2(new_n479), .B1(new_n473), .B2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2067), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n743), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n565), .B2(new_n743), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  NAND3_X1  g348(.A1(new_n760), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT94), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n748), .A2(G2090), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n743), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT23), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n756), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n743), .A2(G24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n613), .B2(new_n743), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1986), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n473), .A2(G131), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n479), .A2(G119), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n478), .A2(G107), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G25), .B(new_n791), .S(G29), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n743), .A2(G23), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n743), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT33), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1976), .ZN(new_n801));
  NAND2_X1  g376(.A1(G166), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G16), .B2(G22), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT91), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n806), .B(new_n808), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n803), .A2(new_n804), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n801), .A2(new_n805), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n796), .B1(new_n812), .B2(KEYINPUT34), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT92), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n812), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT36), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n815), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n783), .B1(new_n818), .B2(new_n820), .ZN(G311));
  INV_X1    g396(.A(new_n783), .ZN(new_n822));
  INV_X1    g397(.A(new_n820), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n819), .B1(new_n815), .B2(new_n816), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(new_n633), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n507), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n561), .A2(new_n833), .B1(new_n536), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n560), .A2(new_n564), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n564), .ZN(new_n837));
  INV_X1    g412(.A(new_n835), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n837), .A2(new_n838), .A3(new_n559), .A4(new_n831), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n827), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  INV_X1    g417(.A(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n832), .A2(new_n835), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n843), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(G145));
  INV_X1    g424(.A(G37), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n768), .B(new_n495), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n724), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(new_n714), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n479), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n478), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G142), .B2(new_n473), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(new_n647), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n791), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n853), .A2(new_n860), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n476), .B(new_n644), .ZN(new_n864));
  XNOR2_X1  g439(.A(G162), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT99), .B1(new_n853), .B2(new_n860), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n861), .B(new_n865), .C1(new_n867), .C2(new_n862), .ZN(new_n868));
  OAI221_X1 g443(.A(new_n850), .B1(new_n863), .B2(new_n865), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g445(.A1(G303), .A2(G305), .ZN(new_n871));
  NAND2_X1  g446(.A1(G303), .A2(G305), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n613), .B(G288), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n573), .A2(new_n619), .A3(new_n623), .A4(new_n579), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n573), .A2(new_n579), .B1(new_n619), .B2(new_n623), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT41), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g459(.A1(G299), .A2(new_n624), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n879), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n882), .A2(KEYINPUT100), .A3(new_n886), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n840), .B(new_n636), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n882), .B(new_n890), .S(new_n891), .Z(new_n892));
  XOR2_X1   g467(.A(new_n878), .B(new_n892), .Z(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G868), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G868), .B2(new_n846), .ZN(G295));
  OAI21_X1  g470(.A(new_n894), .B1(G868), .B2(new_n846), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n545), .A2(new_n547), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n898), .A2(new_n588), .A3(new_n584), .A4(new_n585), .ZN(new_n899));
  NAND2_X1  g474(.A1(G286), .A2(G171), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(G168), .A2(KEYINPUT102), .A3(new_n585), .A4(new_n584), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(new_n840), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n840), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT103), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n840), .A3(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n882), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n883), .A2(new_n887), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n904), .A2(new_n905), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n877), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n901), .B1(new_n586), .B2(G286), .ZN(new_n917));
  AND2_X1   g492(.A1(G286), .A2(G171), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n903), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n840), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n902), .A2(new_n840), .A3(new_n903), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n882), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n882), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n908), .B1(new_n921), .B2(new_n922), .ZN(new_n928));
  INV_X1    g503(.A(new_n909), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n890), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n877), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n915), .A2(new_n916), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n931), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n877), .B1(new_n927), .B2(new_n930), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(G37), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n906), .A2(new_n909), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n937), .A2(new_n890), .B1(new_n925), .B2(new_n926), .ZN(new_n938));
  OAI211_X1 g513(.A(KEYINPUT105), .B(new_n850), .C1(new_n938), .C2(new_n877), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n933), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n897), .B(new_n932), .C1(new_n940), .C2(new_n916), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n931), .A2(new_n916), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n936), .B2(new_n939), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n916), .B1(new_n915), .B2(new_n931), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(G397));
  OR2_X1    g521(.A1(G290), .A2(G1986), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n768), .B(G2067), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n724), .B(G1996), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n791), .B(new_n793), .ZN(new_n951));
  NAND2_X1  g526(.A1(G290), .A2(G1986), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT106), .B(G1384), .Z(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(G164), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n468), .A2(G40), .A3(new_n475), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G1384), .B1(new_n490), .B2(new_n494), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  INV_X1    g538(.A(G1956), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT114), .ZN(new_n966));
  OR3_X1    g541(.A1(G164), .A2(new_n954), .A3(new_n955), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n495), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n957), .B1(new_n969), .B2(new_n954), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(new_n717), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n976));
  AOI21_X1  g551(.A(G299), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n977), .B(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n980), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n957), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n960), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G2067), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n960), .A2(KEYINPUT107), .A3(new_n961), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n962), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT117), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n962), .C1(new_n988), .C2(new_n989), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n986), .B1(new_n994), .B2(new_n759), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n624), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT118), .B(new_n981), .C1(new_n983), .C2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n981), .B1(new_n983), .B2(new_n996), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT61), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n974), .A2(new_n980), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n983), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT61), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT58), .B(G1341), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n985), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n967), .A2(new_n970), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(G1996), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n565), .C1(KEYINPUT119), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(KEYINPUT119), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1003), .A2(new_n1004), .A3(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT120), .B(new_n633), .C1(new_n995), .C2(KEYINPUT60), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n624), .B(KEYINPUT120), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n995), .A2(KEYINPUT60), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n995), .A2(KEYINPUT60), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n997), .B(new_n1000), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT125), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n985), .C1(G288), .C2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(KEYINPUT52), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n985), .A2(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n798), .B2(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1021), .A3(new_n1027), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n601), .A2(new_n605), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n511), .B1(new_n598), .B2(new_n599), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n1034), .B2(new_n604), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT111), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1033), .A2(new_n1035), .A3(new_n1038), .A4(KEYINPUT49), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT49), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n1025), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1040), .A2(KEYINPUT112), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT112), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1031), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT113), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1031), .B(new_n1047), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n969), .A2(new_n954), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n960), .A2(KEYINPUT45), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n984), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1966), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2084), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n962), .C1(new_n988), .C2(new_n989), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1051), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G286), .A2(G8), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1050), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1063), .B(new_n1060), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT121), .B1(new_n1065), .B2(new_n1061), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1062), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(G8), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT51), .A3(new_n1060), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT122), .B(G1961), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n991), .A2(new_n993), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1007), .B2(G2078), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n737), .A2(KEYINPUT123), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n737), .A2(KEYINPUT123), .ZN(new_n1077));
  NOR4_X1   g652(.A1(new_n957), .A2(new_n1074), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n967), .A2(new_n956), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1071), .B1(new_n1080), .B2(G171), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n970), .A2(KEYINPUT53), .A3(new_n737), .A4(new_n1053), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1073), .A2(G301), .A3(new_n1075), .A4(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1068), .A2(new_n1070), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G303), .A2(G8), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1085), .B(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1007), .A2(new_n804), .ZN(new_n1089));
  INV_X1    g664(.A(G2090), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n962), .C1(new_n988), .C2(new_n989), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT108), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(KEYINPUT108), .A3(new_n1091), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1088), .A2(new_n1094), .A3(G8), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1089), .B1(G2090), .B2(new_n963), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G8), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1085), .B(new_n1086), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1049), .A2(new_n1084), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1073), .A2(new_n1075), .A3(new_n1082), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n586), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1073), .A2(G301), .A3(new_n1075), .A4(new_n1079), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1108), .B2(new_n1071), .ZN(new_n1109));
  AOI211_X1 g684(.A(KEYINPUT124), .B(KEYINPUT54), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1020), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT54), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(new_n1104), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1101), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(KEYINPUT125), .A3(new_n1115), .A4(new_n1084), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1019), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1040), .A2(KEYINPUT112), .A3(new_n1042), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1047), .B1(new_n1122), .B2(new_n1031), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1048), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1102), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1070), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT62), .B1(new_n1067), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1106), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1065), .A2(new_n1061), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1063), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1065), .A2(KEYINPUT121), .A3(new_n1061), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1070), .A4(new_n1062), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1127), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT126), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1127), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1115), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1096), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1059), .A2(G168), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1045), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1094), .A2(G8), .A3(new_n1095), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1144), .B(new_n1145), .C1(new_n1088), .C2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1143), .B(new_n1101), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(KEYINPUT63), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1122), .A2(new_n1022), .A3(new_n798), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1025), .B1(new_n1150), .B2(new_n1033), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1145), .B2(new_n1141), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1140), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n959), .B1(new_n1117), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n958), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n791), .A2(new_n794), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n950), .A2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n768), .A2(G2067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OR3_X1    g734(.A1(new_n956), .A2(G1996), .A3(new_n957), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT46), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n958), .B1(new_n724), .B2(new_n948), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT47), .Z(new_n1164));
  NOR2_X1   g739(.A1(new_n947), .A2(new_n1155), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1165), .A2(KEYINPUT48), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1155), .B1(new_n950), .B2(new_n951), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(KEYINPUT48), .B2(new_n1165), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1159), .B(new_n1164), .C1(new_n1166), .C2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT127), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1154), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g746(.A(new_n932), .B1(new_n940), .B2(new_n916), .ZN(new_n1173));
  NOR4_X1   g747(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n1173), .A2(new_n869), .A3(new_n1174), .ZN(G308));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n869), .A3(new_n1174), .ZN(G225));
endmodule


