//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n191), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n193), .B(new_n188), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT65), .B1(new_n200), .B2(G134), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n203), .B2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT66), .A2(G131), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n207), .A2(new_n208), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n210), .A3(new_n205), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n199), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n205), .A2(new_n216), .A3(new_n207), .A4(new_n208), .ZN(new_n217));
  XNOR2_X1  g031(.A(G134), .B(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT67), .B1(new_n218), .B2(new_n216), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n200), .A2(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G131), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(G128), .B(new_n226), .C1(new_n195), .C2(new_n197), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n196), .A2(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n194), .A2(G146), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n228), .B(new_n229), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n215), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n237), .B2(new_n238), .ZN(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n241), .B(new_n243), .C1(new_n237), .C2(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(new_n225), .B2(new_n232), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n235), .A2(KEYINPUT70), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n192), .A2(new_n198), .ZN(new_n251));
  INV_X1    g065(.A(new_n214), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n210), .B1(new_n213), .B2(new_n205), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n223), .B1(new_n222), .B2(G131), .ZN(new_n255));
  AOI211_X1 g069(.A(KEYINPUT67), .B(new_n216), .C1(new_n220), .C2(new_n221), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n227), .A2(new_n231), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n234), .A4(new_n217), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n249), .A2(new_n254), .A3(new_n248), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n262), .A3(KEYINPUT28), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n233), .A2(new_n215), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT28), .B1(new_n264), .B2(new_n248), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n248), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(G237), .A2(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G210), .ZN(new_n270));
  INV_X1    g084(.A(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n187), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  AOI211_X1 g090(.A(KEYINPUT72), .B(new_n274), .C1(new_n263), .C2(new_n267), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n249), .A2(new_n254), .A3(new_n259), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT30), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n264), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n247), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n250), .A2(new_n262), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .A4(new_n274), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(new_n286), .A3(new_n274), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n288), .A3(KEYINPUT31), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n278), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G472), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n279), .A2(new_n247), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n302));
  INV_X1    g116(.A(new_n265), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n275), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n296), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n296), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n283), .A2(new_n247), .B1(new_n250), .B2(new_n262), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(new_n274), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(new_n304), .C1(new_n275), .C2(new_n268), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n295), .A4(new_n296), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n299), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT16), .B1(new_n318), .B2(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT76), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(KEYINPUT76), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n319), .B1(new_n323), .B2(KEYINPUT16), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n324), .A2(new_n196), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n196), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n230), .A2(G119), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G110), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(KEYINPUT75), .A3(G128), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n336), .A2(new_n337), .B1(G119), .B2(new_n230), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT24), .B(G110), .Z(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n325), .B(new_n327), .C1(new_n334), .C2(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n333), .A2(G110), .B1(new_n338), .B2(new_n339), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n324), .A2(new_n196), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n324), .A2(new_n196), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n346), .B(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n349), .B1(new_n341), .B2(new_n345), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G234), .ZN(new_n354));
  OAI21_X1  g168(.A(G217), .B1(new_n354), .B2(G902), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n296), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n355), .B(KEYINPUT74), .Z(new_n359));
  NOR3_X1   g173(.A1(new_n351), .A2(new_n352), .A3(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(KEYINPUT78), .B2(KEYINPUT25), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n341), .A2(new_n345), .ZN(new_n364));
  INV_X1    g178(.A(new_n349), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n296), .A4(new_n350), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT25), .B1(new_n367), .B2(KEYINPUT78), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n358), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G475), .A2(G902), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n343), .A2(new_n344), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n269), .A2(G143), .A3(G214), .ZN(new_n373));
  AOI21_X1  g187(.A(G143), .B1(new_n269), .B2(G214), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n216), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT17), .ZN(new_n377));
  OAI21_X1  g191(.A(G131), .B1(new_n373), .B2(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n372), .B(new_n379), .C1(new_n377), .C2(new_n378), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n323), .A2(G146), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n375), .A2(new_n381), .B1(new_n382), .B2(new_n327), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT18), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n378), .ZN(new_n385));
  XNOR2_X1  g199(.A(G113), .B(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT91), .B(G104), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n380), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n344), .B1(new_n378), .B2(new_n376), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT19), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n393), .B1(new_n321), .B2(new_n322), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT90), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT90), .B1(new_n326), .B2(new_n393), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(new_n394), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(G146), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n389), .B1(new_n399), .B2(new_n385), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n371), .B1(new_n391), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(KEYINPUT20), .B2(new_n401), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n389), .B1(new_n380), .B2(new_n385), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n296), .B1(new_n391), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G475), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G122), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G116), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT92), .ZN(new_n411));
  INV_X1    g225(.A(G116), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G122), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G107), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n411), .B(new_n413), .C1(KEYINPUT14), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n194), .A2(G128), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n230), .A2(G143), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n421), .A2(KEYINPUT93), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(KEYINPUT93), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n203), .ZN(new_n425));
  AOI21_X1  g239(.A(G134), .B1(new_n422), .B2(new_n423), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n416), .B(new_n418), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n203), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n420), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n419), .A2(new_n429), .ZN(new_n432));
  OAI21_X1  g246(.A(G134), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n414), .A2(G107), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n417), .B1(new_n411), .B2(new_n413), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n428), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT9), .B(G234), .Z(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(G217), .A3(new_n347), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n427), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n427), .B2(new_n436), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n296), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n442), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(G234), .A2(G237), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n446), .A2(G952), .A3(new_n347), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT21), .B(G898), .Z(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n446), .A2(G902), .A3(G953), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n408), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G224), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G953), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n456));
  INV_X1    g270(.A(G125), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n192), .B2(new_n198), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  AOI21_X1  g274(.A(G125), .B1(new_n227), .B2(new_n231), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT88), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n456), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT8), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n417), .A2(G104), .ZN(new_n468));
  INV_X1    g282(.A(G104), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G107), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n271), .B1(new_n468), .B2(new_n470), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n417), .A3(G104), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT3), .B1(new_n469), .B2(G107), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n469), .A2(G107), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n271), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n412), .A2(KEYINPUT5), .A3(G119), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n238), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT5), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(new_n244), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n477), .A2(new_n482), .B1(new_n246), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n473), .B(new_n271), .C1(new_n468), .C2(new_n470), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n482), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n246), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n467), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G101), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n497), .A3(G101), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n247), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n477), .A2(new_n246), .A3(new_n482), .A4(new_n486), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n466), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n459), .A2(KEYINPUT7), .A3(new_n463), .A4(new_n455), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n465), .A2(new_n493), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n503), .A2(new_n296), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  INV_X1    g319(.A(new_n466), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n459), .A2(new_n455), .A3(new_n463), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n454), .B1(new_n458), .B2(new_n461), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT87), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT87), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n514), .A3(new_n506), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G210), .B1(G237), .B2(G902), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n504), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n504), .B2(new_n516), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G214), .B1(G237), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n437), .ZN(new_n524));
  OAI21_X1  g338(.A(G221), .B1(new_n524), .B2(G902), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT80), .Z(new_n526));
  INV_X1    g340(.A(G469), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n490), .B2(new_n232), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT10), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT82), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n477), .A2(new_n258), .A3(new_n482), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n252), .A2(new_n253), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n496), .A2(new_n251), .A3(new_n498), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n529), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT83), .B1(new_n212), .B2(new_n214), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n490), .A2(new_n232), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n258), .B1(new_n477), .B2(new_n482), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n536), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  XNOR2_X1  g358(.A(G110), .B(G140), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n347), .A2(G227), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n545), .B(new_n546), .Z(new_n547));
  NAND4_X1  g361(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n529), .A2(new_n534), .A3(new_n532), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(KEYINPUT84), .B2(new_n533), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n533), .A2(KEYINPUT84), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n534), .A3(new_n532), .A4(new_n529), .ZN(new_n552));
  INV_X1    g366(.A(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT86), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n550), .A2(new_n552), .A3(new_n556), .A4(new_n553), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n548), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n544), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n541), .B2(new_n537), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n543), .B1(new_n560), .B2(new_n547), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n527), .B(new_n296), .C1(new_n558), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n550), .A2(new_n552), .A3(new_n547), .ZN(new_n563));
  INV_X1    g377(.A(new_n560), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n547), .ZN(new_n565));
  OAI21_X1  g379(.A(G469), .B1(new_n565), .B2(G902), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n526), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n452), .A2(new_n523), .A3(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n317), .A2(new_n370), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n271), .ZN(G3));
  INV_X1    g384(.A(new_n451), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n521), .B(new_n571), .C1(new_n518), .C2(new_n519), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n567), .A2(new_n370), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n294), .A2(new_n296), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G472), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n574), .A2(new_n297), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n443), .A2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n440), .A2(new_n441), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT33), .B1(new_n441), .B2(KEYINPUT94), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n442), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(G478), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n408), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n577), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT34), .B(G104), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(new_n400), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n390), .ZN(new_n593));
  INV_X1    g407(.A(new_n402), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n371), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n403), .A2(new_n595), .B1(G475), .B2(new_n406), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n596), .A2(new_n445), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n577), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT35), .B(G107), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G9));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n363), .A2(new_n368), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n364), .B1(KEYINPUT36), .B2(new_n365), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n365), .A2(KEYINPUT36), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n341), .A2(new_n345), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n357), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n603), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n608), .B(KEYINPUT97), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(KEYINPUT98), .C1(new_n368), .C2(new_n363), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n567), .A2(new_n523), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n615), .A2(new_n576), .A3(new_n297), .A4(new_n452), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT37), .B(G110), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  AND2_X1   g432(.A1(new_n317), .A2(new_n615), .ZN(new_n619));
  INV_X1    g433(.A(G900), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n447), .B1(new_n450), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n596), .A2(new_n445), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  NAND2_X1  g440(.A1(new_n301), .A2(new_n275), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n628), .A2(new_n290), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n630), .B2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n299), .A2(new_n316), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n520), .B(KEYINPUT38), .Z(new_n633));
  NAND2_X1  g447(.A1(new_n408), .A2(new_n445), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n604), .A2(new_n610), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n634), .A2(new_n636), .A3(new_n522), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT100), .ZN(new_n640));
  INV_X1    g454(.A(new_n567), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n621), .B(KEYINPUT39), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT40), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G143), .ZN(G45));
  NAND2_X1  g460(.A1(new_n588), .A2(new_n622), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n619), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  NOR2_X1   g464(.A1(new_n558), .A2(new_n561), .ZN(new_n651));
  OAI21_X1  g465(.A(G469), .B1(new_n651), .B2(G902), .ZN(new_n652));
  INV_X1    g466(.A(new_n526), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n562), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n587), .A2(new_n572), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n317), .A2(new_n370), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT41), .B(G113), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G15));
  AND2_X1   g473(.A1(new_n597), .A2(new_n573), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n317), .A2(new_n660), .A3(new_n370), .A4(new_n655), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  NAND2_X1  g476(.A1(new_n452), .A2(new_n614), .ZN(new_n663));
  INV_X1    g477(.A(new_n523), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n664), .A3(new_n654), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(new_n317), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n330), .ZN(G21));
  NOR3_X1   g481(.A1(new_n654), .A2(new_n572), .A3(new_n634), .ZN(new_n668));
  NOR2_X1   g482(.A1(G472), .A2(G902), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n291), .A2(new_n287), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n302), .A2(new_n303), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n275), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n575), .B2(G472), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n668), .A2(new_n675), .A3(new_n370), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT101), .B(G122), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G24));
  NOR2_X1   g492(.A1(new_n654), .A2(new_n664), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT102), .B1(new_n675), .B2(new_n636), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n681), .A2(new_n682), .A3(new_n635), .A4(new_n674), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n648), .B(new_n679), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  INV_X1    g499(.A(new_n519), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n504), .A2(new_n516), .A3(new_n517), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n521), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n641), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n317), .A2(new_n691), .A3(new_n370), .A4(new_n648), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT104), .B(G131), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G33));
  XOR2_X1   g510(.A(new_n623), .B(KEYINPUT105), .Z(new_n697));
  NAND4_X1  g511(.A1(new_n317), .A2(new_n691), .A3(new_n370), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G134), .ZN(G36));
  OR2_X1    g513(.A1(new_n565), .A2(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n565), .A2(KEYINPUT45), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(G469), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(G469), .A2(G902), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n562), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n653), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(new_n642), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n690), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n576), .A2(new_n297), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n636), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT107), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n584), .A2(new_n586), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n408), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT43), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n713), .A2(new_n714), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G137), .ZN(G39));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n710), .A2(new_n728), .A3(new_n653), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n710), .B2(new_n653), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n648), .A2(new_n369), .A3(new_n714), .ZN(new_n732));
  OR4_X1    g546(.A1(new_n317), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G140), .ZN(G42));
  OR2_X1    g548(.A1(new_n632), .A2(new_n369), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n652), .A2(new_n562), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(KEYINPUT49), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(KEYINPUT49), .ZN(new_n738));
  INV_X1    g552(.A(new_n633), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n521), .A3(new_n653), .A4(new_n720), .ZN(new_n740));
  OR4_X1    g554(.A1(new_n735), .A2(new_n737), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n744));
  INV_X1    g558(.A(new_n674), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n576), .A2(new_n745), .A3(new_n636), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n682), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n675), .A2(KEYINPUT102), .A3(new_n636), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT109), .A3(new_n648), .A4(new_n691), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n648), .B(new_n691), .C1(new_n680), .C2(new_n683), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n596), .A2(new_n622), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n445), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n444), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n585), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n442), .A2(new_n444), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT108), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n755), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n317), .A2(new_n614), .A3(new_n691), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n698), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n744), .B1(new_n754), .B2(new_n765), .ZN(new_n766));
  AOI211_X1 g580(.A(KEYINPUT110), .B(new_n764), .C1(new_n750), .C2(new_n753), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n317), .B(new_n615), .C1(new_n624), .C2(new_n648), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n684), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n635), .A2(new_n622), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n641), .A2(new_n664), .A3(new_n634), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n632), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n774), .B1(new_n632), .B2(new_n773), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n769), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n632), .A2(new_n773), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n632), .A2(new_n773), .A3(new_n774), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(KEYINPUT52), .A3(new_n684), .A4(new_n770), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n657), .A2(new_n661), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n404), .A2(new_n407), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n757), .B2(new_n761), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n587), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n574), .A2(new_n788), .A3(new_n297), .A4(new_n576), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n676), .A2(new_n616), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n666), .ZN(new_n791));
  INV_X1    g605(.A(new_n569), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n692), .B(KEYINPUT42), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n743), .B1(new_n768), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n751), .A2(new_n752), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n751), .A2(new_n752), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n765), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT110), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n754), .A2(new_n744), .A3(new_n765), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n790), .A2(new_n569), .A3(new_n666), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n694), .A2(new_n805), .A3(new_n785), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n778), .B2(new_n783), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n804), .A2(new_n807), .A3(KEYINPUT53), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n797), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n798), .B1(new_n797), .B2(new_n808), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n742), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n768), .A2(new_n796), .A3(new_n743), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT53), .B1(new_n804), .B2(new_n807), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT54), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n797), .A2(new_n808), .A3(new_n798), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(KEYINPUT112), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n721), .A2(new_n447), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n818), .A2(new_n370), .A3(new_n675), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n522), .A2(new_n819), .A3(new_n739), .A4(new_n655), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT50), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n714), .A2(KEYINPUT113), .A3(new_n655), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n690), .B2(new_n654), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n447), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n735), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n408), .A2(new_n584), .A3(new_n586), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n821), .A2(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n730), .A2(new_n731), .B1(new_n653), .B2(new_n736), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n819), .A2(new_n714), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n818), .A2(new_n825), .A3(new_n823), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT114), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n830), .A2(new_n831), .B1(new_n749), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n829), .B2(new_n834), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n819), .A2(new_n523), .A3(new_n655), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(G952), .A3(new_n347), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n588), .B2(new_n827), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT48), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n317), .A2(new_n370), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n833), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n840), .B1(new_n833), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n835), .A2(new_n836), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n817), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(G952), .B2(G953), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n817), .B2(new_n845), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n741), .B1(new_n848), .B2(new_n849), .ZN(G75));
  NOR2_X1   g664(.A1(new_n347), .A2(G952), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n797), .A2(new_n808), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(G210), .A3(G902), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n508), .A2(new_n515), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(new_n513), .Z(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT55), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n852), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT56), .B1(new_n854), .B2(KEYINPUT116), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(KEYINPUT116), .B2(new_n854), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n858), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(KEYINPUT117), .A3(new_n858), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(G51));
  AOI21_X1  g681(.A(new_n296), .B1(new_n797), .B2(new_n808), .ZN(new_n868));
  INV_X1    g682(.A(new_n702), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n814), .A2(new_n815), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n703), .B(KEYINPUT57), .Z(new_n874));
  AOI21_X1  g688(.A(new_n651), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n852), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n878), .B(new_n852), .C1(new_n872), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  INV_X1    g695(.A(new_n593), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n851), .ZN(G60));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  NAND2_X1  g700(.A1(G478), .A2(G902), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT59), .Z(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n811), .A2(new_n816), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n582), .A2(new_n583), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n888), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n809), .B2(new_n810), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n851), .B1(new_n895), .B2(KEYINPUT120), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n873), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n886), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n890), .A2(new_n892), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n898), .A4(new_n896), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(G63));
  OAI21_X1  g717(.A(new_n852), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT60), .Z(new_n906));
  AND2_X1   g720(.A1(new_n853), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n353), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n605), .A2(new_n607), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(KEYINPUT122), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n907), .B2(new_n912), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n910), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n907), .A2(new_n912), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n913), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n911), .B1(new_n921), .B2(new_n910), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n917), .A2(new_n922), .ZN(G66));
  OAI21_X1  g737(.A(G953), .B1(new_n449), .B2(new_n453), .ZN(new_n924));
  INV_X1    g738(.A(new_n793), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n856), .B1(G898), .B2(new_n347), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT124), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  INV_X1    g743(.A(new_n698), .ZN(new_n930));
  INV_X1    g744(.A(new_n841), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n931), .A2(new_n664), .A3(new_n634), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n794), .B(new_n930), .C1(new_n713), .C2(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n771), .B(KEYINPUT125), .Z(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n726), .A3(new_n733), .A4(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n283), .B(new_n398), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(G900), .B2(G953), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n733), .A2(new_n726), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n841), .A2(new_n691), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n788), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n642), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n934), .A2(new_n645), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  AOI21_X1  g763(.A(G953), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n937), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n939), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n347), .B1(G227), .B2(G900), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n939), .B(new_n955), .C1(new_n950), .C2(new_n951), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G72));
  NAND3_X1  g771(.A1(new_n947), .A2(new_n925), .A3(new_n949), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n959));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n275), .B(new_n311), .C1(new_n958), .C2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n935), .B2(new_n793), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n963), .A2(new_n275), .A3(new_n311), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n312), .A2(new_n290), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n853), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n962), .A2(new_n851), .A3(new_n964), .A4(new_n966), .ZN(G57));
endmodule


