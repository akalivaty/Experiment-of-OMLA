

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734;

  NOR2_X1 U366 ( .A1(n697), .A2(n706), .ZN(n364) );
  NOR2_X1 U367 ( .A1(n620), .A2(n706), .ZN(n621) );
  AND2_X1 U368 ( .A1(n384), .A2(n387), .ZN(n383) );
  XNOR2_X1 U369 ( .A(n524), .B(n422), .ZN(n729) );
  XNOR2_X1 U370 ( .A(n492), .B(KEYINPUT39), .ZN(n567) );
  NOR2_X1 U371 ( .A1(n629), .A2(n630), .ZN(n593) );
  NOR2_X1 U372 ( .A1(n553), .A2(n630), .ZN(n597) );
  NAND2_X1 U373 ( .A1(n347), .A2(n346), .ZN(n399) );
  XNOR2_X1 U374 ( .A(n592), .B(n348), .ZN(n347) );
  INV_X1 U375 ( .A(n354), .ZN(n346) );
  INV_X1 U376 ( .A(n476), .ZN(n348) );
  XNOR2_X1 U377 ( .A(n345), .B(n344), .ZN(n472) );
  XNOR2_X1 U378 ( .A(n469), .B(n468), .ZN(n344) );
  INV_X1 U379 ( .A(KEYINPUT65), .ZN(n369) );
  NAND2_X2 U380 ( .A1(n343), .A2(n375), .ZN(n700) );
  NAND2_X1 U381 ( .A1(n606), .A2(n373), .ZN(n343) );
  XNOR2_X2 U382 ( .A(n508), .B(G134), .ZN(n368) );
  INV_X1 U383 ( .A(n484), .ZN(n345) );
  XOR2_X1 U384 ( .A(G137), .B(G140), .Z(n452) );
  XNOR2_X1 U385 ( .A(n553), .B(KEYINPUT1), .ZN(n629) );
  NOR2_X1 U386 ( .A1(n609), .A2(G902), .ZN(n475) );
  XNOR2_X1 U387 ( .A(n474), .B(n473), .ZN(n609) );
  AND2_X2 U388 ( .A1(n427), .A2(n365), .ZN(n605) );
  NAND2_X1 U389 ( .A1(n623), .A2(n622), .ZN(n630) );
  NOR2_X1 U390 ( .A1(n603), .A2(n579), .ZN(n581) );
  XNOR2_X1 U391 ( .A(n496), .B(n485), .ZN(n486) );
  NOR2_X1 U392 ( .A1(n612), .A2(n706), .ZN(n615) );
  OR2_X1 U393 ( .A1(n563), .A2(n386), .ZN(n382) );
  NOR2_X1 U394 ( .A1(n412), .A2(n411), .ZN(n410) );
  NAND2_X1 U395 ( .A1(n562), .A2(n388), .ZN(n387) );
  XNOR2_X1 U396 ( .A(n581), .B(n580), .ZN(n732) );
  NAND2_X1 U397 ( .A1(n380), .A2(n352), .ZN(n379) );
  XNOR2_X1 U398 ( .A(n403), .B(n402), .ZN(n730) );
  XNOR2_X1 U399 ( .A(n430), .B(n381), .ZN(n380) );
  NOR2_X1 U400 ( .A1(n396), .A2(n395), .ZN(n477) );
  OR2_X1 U401 ( .A1(n702), .A2(G902), .ZN(n433) );
  XNOR2_X1 U402 ( .A(n467), .B(G113), .ZN(n484) );
  XNOR2_X1 U403 ( .A(G101), .B(KEYINPUT3), .ZN(n467) );
  XNOR2_X1 U404 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n370) );
  BUF_X1 U405 ( .A(n700), .Z(n349) );
  XNOR2_X1 U406 ( .A(n592), .B(n476), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X2 U408 ( .A(n368), .B(n482), .ZN(n716) );
  XNOR2_X2 U409 ( .A(n716), .B(G146), .ZN(n474) );
  XNOR2_X1 U410 ( .A(n418), .B(G146), .ZN(n480) );
  INV_X1 U411 ( .A(G125), .ZN(n418) );
  NAND2_X1 U412 ( .A1(n672), .A2(n585), .ZN(n408) );
  OR2_X1 U413 ( .A1(n732), .A2(n406), .ZN(n405) );
  INV_X1 U414 ( .A(n585), .ZN(n406) );
  XNOR2_X1 U415 ( .A(n451), .B(KEYINPUT10), .ZN(n506) );
  OR2_X1 U416 ( .A1(G902), .A2(G237), .ZN(n490) );
  XNOR2_X1 U417 ( .A(n414), .B(KEYINPUT0), .ZN(n591) );
  NOR2_X1 U418 ( .A1(n575), .A2(n574), .ZN(n414) );
  INV_X1 U419 ( .A(KEYINPUT78), .ZN(n420) );
  XNOR2_X1 U420 ( .A(n498), .B(n361), .ZN(n502) );
  AND2_X1 U421 ( .A1(n600), .A2(n366), .ZN(n365) );
  NOR2_X1 U422 ( .A1(n548), .A2(n730), .ZN(n549) );
  AND2_X1 U423 ( .A1(G953), .A2(G902), .ZN(n463) );
  XOR2_X1 U424 ( .A(G134), .B(KEYINPUT92), .Z(n494) );
  NOR2_X1 U425 ( .A1(G953), .A2(G237), .ZN(n505) );
  INV_X1 U426 ( .A(KEYINPUT72), .ZN(n416) );
  XNOR2_X1 U427 ( .A(n480), .B(n481), .ZN(n417) );
  OR2_X1 U428 ( .A1(n731), .A2(KEYINPUT44), .ZN(n428) );
  XOR2_X1 U429 ( .A(KEYINPUT71), .B(KEYINPUT23), .Z(n448) );
  XNOR2_X1 U430 ( .A(G128), .B(KEYINPUT24), .ZN(n447) );
  XNOR2_X1 U431 ( .A(n511), .B(n367), .ZN(n694) );
  XNOR2_X1 U432 ( .A(n517), .B(n510), .ZN(n367) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n510) );
  XNOR2_X1 U434 ( .A(n589), .B(KEYINPUT101), .ZN(n431) );
  INV_X1 U435 ( .A(KEYINPUT33), .ZN(n589) );
  NOR2_X1 U436 ( .A1(n553), .A2(n531), .ZN(n539) );
  XNOR2_X1 U437 ( .A(n530), .B(n529), .ZN(n531) );
  INV_X1 U438 ( .A(n550), .ZN(n362) );
  XNOR2_X1 U439 ( .A(n504), .B(KEYINPUT94), .ZN(n545) );
  XNOR2_X1 U440 ( .A(n413), .B(n358), .ZN(n582) );
  NAND2_X1 U441 ( .A1(n576), .A2(n591), .ZN(n413) );
  AND2_X1 U442 ( .A1(n642), .A2(n622), .ZN(n576) );
  XNOR2_X1 U443 ( .A(n458), .B(n353), .ZN(n432) );
  NAND2_X1 U444 ( .A1(n378), .A2(n376), .ZN(n375) );
  NOR2_X1 U445 ( .A1(n608), .A2(n377), .ZN(n376) );
  XNOR2_X1 U446 ( .A(n426), .B(n423), .ZN(n438) );
  NOR2_X1 U447 ( .A1(G952), .A2(n443), .ZN(n706) );
  INV_X1 U448 ( .A(KEYINPUT48), .ZN(n388) );
  NAND2_X1 U449 ( .A1(G237), .A2(G234), .ZN(n461) );
  NOR2_X1 U450 ( .A1(n672), .A2(n585), .ZN(n411) );
  XNOR2_X1 U451 ( .A(n499), .B(n355), .ZN(n361) );
  XNOR2_X1 U452 ( .A(G122), .B(KEYINPUT9), .ZN(n493) );
  XNOR2_X1 U453 ( .A(n506), .B(n507), .ZN(n509) );
  INV_X1 U454 ( .A(n666), .ZN(n366) );
  INV_X1 U455 ( .A(KEYINPUT28), .ZN(n528) );
  XOR2_X1 U456 ( .A(KEYINPUT38), .B(n546), .Z(n640) );
  AND2_X1 U457 ( .A1(n400), .A2(n398), .ZN(n397) );
  NAND2_X1 U458 ( .A1(n401), .A2(KEYINPUT30), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n538), .B(KEYINPUT19), .ZN(n570) );
  XNOR2_X1 U460 ( .A(KEYINPUT97), .B(n532), .ZN(n642) );
  XNOR2_X1 U461 ( .A(G122), .B(G104), .ZN(n512) );
  XNOR2_X1 U462 ( .A(G902), .B(KEYINPUT15), .ZN(n608) );
  AND2_X1 U463 ( .A1(n709), .A2(n374), .ZN(n373) );
  INV_X1 U464 ( .A(n608), .ZN(n374) );
  XNOR2_X1 U465 ( .A(n452), .B(n437), .ZN(n426) );
  XNOR2_X1 U466 ( .A(n425), .B(n424), .ZN(n423) );
  XNOR2_X1 U467 ( .A(G101), .B(G110), .ZN(n425) );
  XNOR2_X1 U468 ( .A(G107), .B(G104), .ZN(n424) );
  XNOR2_X1 U469 ( .A(n417), .B(n415), .ZN(n483) );
  XNOR2_X1 U470 ( .A(n479), .B(n416), .ZN(n415) );
  INV_X1 U471 ( .A(KEYINPUT34), .ZN(n381) );
  XNOR2_X1 U472 ( .A(n521), .B(n520), .ZN(n541) );
  XNOR2_X1 U473 ( .A(n453), .B(n717), .ZN(n702) );
  XNOR2_X1 U474 ( .A(n394), .B(n393), .ZN(n392) );
  NAND2_X1 U475 ( .A1(n700), .A2(G478), .ZN(n394) );
  NAND2_X1 U476 ( .A1(n378), .A2(KEYINPUT2), .ZN(n372) );
  XNOR2_X1 U477 ( .A(n536), .B(n535), .ZN(n733) );
  NOR2_X1 U478 ( .A1(n555), .A2(n601), .ZN(n686) );
  INV_X1 U479 ( .A(KEYINPUT32), .ZN(n580) );
  XNOR2_X1 U480 ( .A(KEYINPUT95), .B(n522), .ZN(n676) );
  NAND2_X1 U481 ( .A1(n545), .A2(n541), .ZN(n522) );
  INV_X1 U482 ( .A(KEYINPUT103), .ZN(n402) );
  AND2_X1 U483 ( .A1(n547), .A2(n404), .ZN(n403) );
  AND2_X1 U484 ( .A1(n590), .A2(n546), .ZN(n404) );
  XNOR2_X1 U485 ( .A(n390), .B(n389), .ZN(G63) );
  INV_X1 U486 ( .A(KEYINPUT122), .ZN(n389) );
  NAND2_X1 U487 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U488 ( .A(n706), .ZN(n391) );
  XNOR2_X1 U489 ( .A(n690), .B(n360), .ZN(n692) );
  XNOR2_X1 U490 ( .A(n419), .B(n691), .ZN(n360) );
  AND2_X1 U491 ( .A1(n676), .A2(n357), .ZN(n351) );
  XNOR2_X1 U492 ( .A(n590), .B(KEYINPUT74), .ZN(n352) );
  XOR2_X1 U493 ( .A(n455), .B(n454), .Z(n353) );
  OR2_X1 U494 ( .A1(n401), .A2(KEYINPUT30), .ZN(n354) );
  XOR2_X1 U495 ( .A(KEYINPUT7), .B(KEYINPUT93), .Z(n355) );
  AND2_X1 U496 ( .A1(n372), .A2(n371), .ZN(n356) );
  AND2_X1 U497 ( .A1(n586), .A2(n362), .ZN(n357) );
  XOR2_X1 U498 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n358) );
  XNOR2_X1 U499 ( .A(KEYINPUT73), .B(KEYINPUT35), .ZN(n359) );
  NOR2_X1 U500 ( .A1(n686), .A2(n556), .ZN(n557) );
  XNOR2_X1 U501 ( .A(n489), .B(n712), .ZN(n616) );
  XNOR2_X2 U502 ( .A(n534), .B(KEYINPUT41), .ZN(n656) );
  XNOR2_X1 U503 ( .A(n364), .B(n698), .ZN(G60) );
  XNOR2_X2 U504 ( .A(n369), .B(G131), .ZN(n508) );
  XNOR2_X2 U505 ( .A(n495), .B(n370), .ZN(n482) );
  XNOR2_X2 U506 ( .A(G143), .B(G128), .ZN(n495) );
  NAND2_X1 U507 ( .A1(n709), .A2(n607), .ZN(n378) );
  XNOR2_X2 U508 ( .A(n605), .B(n604), .ZN(n709) );
  NAND2_X1 U509 ( .A1(n606), .A2(n709), .ZN(n371) );
  INV_X1 U510 ( .A(KEYINPUT2), .ZN(n377) );
  INV_X1 U511 ( .A(n731), .ZN(n412) );
  XNOR2_X2 U512 ( .A(n379), .B(n359), .ZN(n731) );
  NAND2_X1 U513 ( .A1(n383), .A2(n382), .ZN(n385) );
  NAND2_X1 U514 ( .A1(n563), .A2(n388), .ZN(n384) );
  XNOR2_X2 U515 ( .A(n607), .B(n420), .ZN(n720) );
  AND2_X2 U516 ( .A1(n385), .A2(n569), .ZN(n607) );
  OR2_X1 U517 ( .A1(n562), .A2(n388), .ZN(n386) );
  INV_X1 U518 ( .A(n699), .ZN(n393) );
  AND2_X1 U519 ( .A1(n350), .A2(KEYINPUT30), .ZN(n395) );
  NAND2_X1 U520 ( .A1(n399), .A2(n397), .ZN(n396) );
  INV_X1 U521 ( .A(n525), .ZN(n400) );
  INV_X1 U522 ( .A(n639), .ZN(n401) );
  NOR2_X2 U523 ( .A1(n720), .A2(KEYINPUT2), .ZN(n606) );
  XNOR2_X2 U524 ( .A(n442), .B(n441), .ZN(n553) );
  NAND2_X1 U525 ( .A1(n655), .A2(n591), .ZN(n430) );
  NAND2_X1 U526 ( .A1(n407), .A2(n405), .ZN(n409) );
  NAND2_X1 U527 ( .A1(n408), .A2(n732), .ZN(n407) );
  NAND2_X1 U528 ( .A1(n410), .A2(n409), .ZN(n429) );
  NOR2_X1 U529 ( .A1(n419), .A2(G902), .ZN(n442) );
  XNOR2_X1 U530 ( .A(n440), .B(n439), .ZN(n419) );
  XNOR2_X1 U531 ( .A(n421), .B(n537), .ZN(n558) );
  NAND2_X1 U532 ( .A1(n733), .A2(n729), .ZN(n421) );
  XNOR2_X1 U533 ( .A(n523), .B(KEYINPUT106), .ZN(n422) );
  NAND2_X1 U534 ( .A1(n429), .A2(n428), .ZN(n427) );
  XNOR2_X2 U535 ( .A(n588), .B(n431), .ZN(n655) );
  XNOR2_X2 U536 ( .A(n433), .B(n432), .ZN(n623) );
  XNOR2_X1 U537 ( .A(n702), .B(n701), .ZN(n703) );
  INV_X1 U538 ( .A(n495), .ZN(n497) );
  XOR2_X1 U539 ( .A(n515), .B(n514), .Z(n434) );
  AND2_X1 U540 ( .A1(G210), .A2(n490), .ZN(n435) );
  XOR2_X1 U541 ( .A(n618), .B(n617), .Z(n436) );
  XNOR2_X1 U542 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n479) );
  INV_X1 U543 ( .A(n688), .ZN(n568) );
  NOR2_X1 U544 ( .A1(n689), .A2(n568), .ZN(n569) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n489) );
  INV_X1 U546 ( .A(KEYINPUT70), .ZN(n454) );
  XNOR2_X1 U547 ( .A(n516), .B(n434), .ZN(n517) );
  XNOR2_X1 U548 ( .A(n528), .B(KEYINPUT104), .ZN(n529) );
  INV_X1 U549 ( .A(KEYINPUT63), .ZN(n613) );
  XNOR2_X1 U550 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U551 ( .A(n613), .B(KEYINPUT82), .ZN(n614) );
  XNOR2_X1 U552 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U553 ( .A(n665), .B(n664), .ZN(G75) );
  INV_X2 U554 ( .A(G953), .ZN(n443) );
  XNOR2_X1 U555 ( .A(n474), .B(KEYINPUT84), .ZN(n440) );
  NAND2_X1 U556 ( .A1(G227), .A2(n443), .ZN(n437) );
  XOR2_X1 U557 ( .A(n438), .B(KEYINPUT85), .Z(n439) );
  XNOR2_X1 U558 ( .A(KEYINPUT66), .B(G469), .ZN(n441) );
  XOR2_X2 U559 ( .A(G119), .B(G110), .Z(n485) );
  XOR2_X1 U560 ( .A(n485), .B(KEYINPUT67), .Z(n446) );
  NAND2_X1 U561 ( .A1(G234), .A2(n443), .ZN(n444) );
  XOR2_X1 U562 ( .A(KEYINPUT8), .B(n444), .Z(n500) );
  NAND2_X1 U563 ( .A1(G221), .A2(n500), .ZN(n445) );
  XNOR2_X1 U564 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U565 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U566 ( .A(n450), .B(n449), .ZN(n453) );
  INV_X1 U567 ( .A(n480), .ZN(n451) );
  XNOR2_X1 U568 ( .A(n452), .B(n506), .ZN(n717) );
  XNOR2_X1 U569 ( .A(KEYINPUT25), .B(KEYINPUT87), .ZN(n455) );
  NAND2_X1 U570 ( .A1(n608), .A2(G234), .ZN(n457) );
  XNOR2_X1 U571 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n457), .B(n456), .ZN(n459) );
  NAND2_X1 U573 ( .A1(G217), .A2(n459), .ZN(n458) );
  NAND2_X1 U574 ( .A1(n459), .A2(G221), .ZN(n460) );
  XOR2_X1 U575 ( .A(KEYINPUT21), .B(n460), .Z(n622) );
  XNOR2_X1 U576 ( .A(n461), .B(KEYINPUT14), .ZN(n464) );
  NAND2_X1 U577 ( .A1(G952), .A2(n464), .ZN(n653) );
  NOR2_X1 U578 ( .A1(G953), .A2(n653), .ZN(n462) );
  XOR2_X1 U579 ( .A(KEYINPUT83), .B(n462), .Z(n573) );
  NAND2_X1 U580 ( .A1(n464), .A2(n463), .ZN(n571) );
  XNOR2_X1 U581 ( .A(KEYINPUT102), .B(n571), .ZN(n465) );
  NOR2_X1 U582 ( .A1(G900), .A2(n465), .ZN(n466) );
  NOR2_X1 U583 ( .A1(n573), .A2(n466), .ZN(n525) );
  XOR2_X1 U584 ( .A(KEYINPUT5), .B(G137), .Z(n469) );
  XNOR2_X1 U585 ( .A(G116), .B(G119), .ZN(n468) );
  NAND2_X1 U586 ( .A1(n505), .A2(G210), .ZN(n471) );
  XNOR2_X2 U587 ( .A(n475), .B(G472), .ZN(n592) );
  INV_X1 U588 ( .A(KEYINPUT99), .ZN(n476) );
  NAND2_X1 U589 ( .A1(G214), .A2(n490), .ZN(n639) );
  NAND2_X1 U590 ( .A1(n597), .A2(n477), .ZN(n478) );
  XNOR2_X1 U591 ( .A(n478), .B(KEYINPUT69), .ZN(n547) );
  NAND2_X1 U592 ( .A1(G224), .A2(n443), .ZN(n481) );
  XOR2_X1 U593 ( .A(KEYINPUT16), .B(n484), .Z(n488) );
  XOR2_X2 U594 ( .A(G116), .B(G107), .Z(n496) );
  XNOR2_X1 U595 ( .A(n486), .B(n512), .ZN(n487) );
  XNOR2_X1 U596 ( .A(n488), .B(n487), .ZN(n712) );
  NAND2_X1 U597 ( .A1(n616), .A2(n608), .ZN(n491) );
  XNOR2_X2 U598 ( .A(n491), .B(n435), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n547), .A2(n640), .ZN(n492) );
  XNOR2_X1 U600 ( .A(n494), .B(n493), .ZN(n499) );
  XOR2_X1 U601 ( .A(n497), .B(n496), .Z(n498) );
  NAND2_X1 U602 ( .A1(G217), .A2(n500), .ZN(n501) );
  XNOR2_X1 U603 ( .A(n502), .B(n501), .ZN(n699) );
  NOR2_X1 U604 ( .A1(n699), .A2(G902), .ZN(n503) );
  XNOR2_X1 U605 ( .A(G478), .B(n503), .ZN(n504) );
  NAND2_X1 U606 ( .A1(n505), .A2(G214), .ZN(n507) );
  XOR2_X1 U607 ( .A(n508), .B(n509), .Z(n511) );
  INV_X1 U608 ( .A(n512), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n513), .B(KEYINPUT11), .ZN(n516) );
  XOR2_X1 U610 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n515) );
  XNOR2_X1 U611 ( .A(G140), .B(KEYINPUT12), .ZN(n514) );
  NOR2_X1 U612 ( .A1(n694), .A2(G902), .ZN(n521) );
  XOR2_X1 U613 ( .A(KEYINPUT91), .B(KEYINPUT13), .Z(n519) );
  XNOR2_X1 U614 ( .A(KEYINPUT90), .B(G475), .ZN(n518) );
  XNOR2_X1 U615 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U616 ( .A1(n567), .A2(n676), .ZN(n524) );
  XOR2_X1 U617 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n523) );
  NOR2_X1 U618 ( .A1(n623), .A2(n525), .ZN(n526) );
  NAND2_X1 U619 ( .A1(n526), .A2(n622), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n550), .A2(n350), .ZN(n530) );
  INV_X1 U621 ( .A(n541), .ZN(n544) );
  NAND2_X1 U622 ( .A1(n545), .A2(n544), .ZN(n532) );
  NAND2_X1 U623 ( .A1(n640), .A2(n639), .ZN(n533) );
  XNOR2_X1 U624 ( .A(KEYINPUT107), .B(n533), .ZN(n645) );
  NAND2_X1 U625 ( .A1(n642), .A2(n645), .ZN(n534) );
  NAND2_X1 U626 ( .A1(n539), .A2(n656), .ZN(n536) );
  XNOR2_X1 U627 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n535) );
  XOR2_X1 U628 ( .A(KEYINPUT46), .B(KEYINPUT80), .Z(n537) );
  NAND2_X1 U629 ( .A1(n546), .A2(n639), .ZN(n538) );
  NAND2_X1 U630 ( .A1(n539), .A2(n570), .ZN(n559) );
  NAND2_X1 U631 ( .A1(n559), .A2(KEYINPUT47), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n540), .B(KEYINPUT76), .ZN(n543) );
  NOR2_X1 U633 ( .A1(n545), .A2(n541), .ZN(n673) );
  NOR2_X1 U634 ( .A1(n676), .A2(n673), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n560), .A2(KEYINPUT47), .ZN(n542) );
  NAND2_X1 U636 ( .A1(n543), .A2(n542), .ZN(n548) );
  NOR2_X1 U637 ( .A1(n545), .A2(n544), .ZN(n590) );
  XNOR2_X1 U638 ( .A(KEYINPUT75), .B(n549), .ZN(n556) );
  XOR2_X1 U639 ( .A(KEYINPUT109), .B(KEYINPUT36), .Z(n552) );
  XOR2_X1 U640 ( .A(KEYINPUT6), .B(n592), .Z(n577) );
  INV_X1 U641 ( .A(n577), .ZN(n586) );
  AND2_X1 U642 ( .A1(n351), .A2(n639), .ZN(n564) );
  NAND2_X1 U643 ( .A1(n564), .A2(n546), .ZN(n551) );
  XNOR2_X1 U644 ( .A(n552), .B(n551), .ZN(n555) );
  INV_X1 U645 ( .A(n629), .ZN(n554) );
  INV_X1 U646 ( .A(n554), .ZN(n601) );
  NAND2_X1 U647 ( .A1(n558), .A2(n557), .ZN(n563) );
  INV_X1 U648 ( .A(n559), .ZN(n677) );
  INV_X1 U649 ( .A(n560), .ZN(n644) );
  NAND2_X1 U650 ( .A1(n677), .A2(n644), .ZN(n561) );
  NOR2_X1 U651 ( .A1(KEYINPUT47), .A2(n561), .ZN(n562) );
  AND2_X1 U652 ( .A1(n601), .A2(n564), .ZN(n565) );
  XNOR2_X1 U653 ( .A(n565), .B(KEYINPUT43), .ZN(n566) );
  NOR2_X1 U654 ( .A1(n546), .A2(n566), .ZN(n689) );
  NAND2_X1 U655 ( .A1(n567), .A2(n673), .ZN(n688) );
  INV_X1 U656 ( .A(n570), .ZN(n575) );
  NOR2_X1 U657 ( .A1(G898), .A2(n571), .ZN(n572) );
  NOR2_X1 U658 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U659 ( .A1(n582), .A2(n577), .ZN(n603) );
  NOR2_X1 U660 ( .A1(n623), .A2(n601), .ZN(n578) );
  XOR2_X1 U661 ( .A(KEYINPUT98), .B(n578), .Z(n579) );
  NAND2_X1 U662 ( .A1(n582), .A2(n350), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n623), .A2(n583), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n584), .A2(n601), .ZN(n672) );
  NOR2_X1 U665 ( .A1(KEYINPUT44), .A2(KEYINPUT81), .ZN(n585) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT100), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U668 ( .A(n591), .ZN(n595) );
  INV_X1 U669 ( .A(n592), .ZN(n627) );
  NAND2_X1 U670 ( .A1(n627), .A2(n593), .ZN(n636) );
  NOR2_X1 U671 ( .A1(n595), .A2(n636), .ZN(n594) );
  XNOR2_X1 U672 ( .A(KEYINPUT31), .B(n594), .ZN(n682) );
  NOR2_X1 U673 ( .A1(n627), .A2(n595), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n668) );
  NAND2_X1 U675 ( .A1(n682), .A2(n668), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n598), .A2(n644), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n599), .B(KEYINPUT96), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n623), .A2(n601), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n666) );
  XNOR2_X1 U680 ( .A(KEYINPUT79), .B(KEYINPUT45), .ZN(n604) );
  NAND2_X1 U681 ( .A1(G472), .A2(n700), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT62), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(G57) );
  NAND2_X1 U685 ( .A1(n700), .A2(G210), .ZN(n619) );
  XNOR2_X1 U686 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT119), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n619), .B(n436), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n621), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U690 ( .A(n356), .B(KEYINPUT77), .Z(n662) );
  NOR2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U692 ( .A(KEYINPUT49), .B(n624), .Z(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(KEYINPUT112), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U695 ( .A(KEYINPUT113), .B(n628), .Z(n634) );
  NAND2_X1 U696 ( .A1(n630), .A2(n601), .ZN(n631) );
  XNOR2_X1 U697 ( .A(n631), .B(KEYINPUT114), .ZN(n632) );
  XNOR2_X1 U698 ( .A(KEYINPUT50), .B(n632), .ZN(n633) );
  NAND2_X1 U699 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U700 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U701 ( .A(KEYINPUT51), .B(n637), .Z(n638) );
  NAND2_X1 U702 ( .A1(n656), .A2(n638), .ZN(n650) );
  NOR2_X1 U703 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U704 ( .A(KEYINPUT115), .B(n641), .ZN(n643) );
  NAND2_X1 U705 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U706 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U707 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U708 ( .A1(n655), .A2(n648), .ZN(n649) );
  NAND2_X1 U709 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U710 ( .A(KEYINPUT52), .B(n651), .Z(n652) );
  NOR2_X1 U711 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U712 ( .A(KEYINPUT116), .B(n654), .Z(n658) );
  NAND2_X1 U713 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U714 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U715 ( .A(KEYINPUT117), .B(n659), .Z(n660) );
  NOR2_X1 U716 ( .A1(G953), .A2(n660), .ZN(n661) );
  NAND2_X1 U717 ( .A1(n662), .A2(n661), .ZN(n665) );
  INV_X1 U718 ( .A(KEYINPUT118), .ZN(n663) );
  XNOR2_X1 U719 ( .A(n663), .B(KEYINPUT53), .ZN(n664) );
  XOR2_X1 U720 ( .A(G101), .B(n666), .Z(G3) );
  INV_X1 U721 ( .A(n676), .ZN(n680) );
  NOR2_X1 U722 ( .A1(n680), .A2(n668), .ZN(n667) );
  XOR2_X1 U723 ( .A(G104), .B(n667), .Z(G6) );
  INV_X1 U724 ( .A(n673), .ZN(n683) );
  NOR2_X1 U725 ( .A1(n683), .A2(n668), .ZN(n670) );
  XNOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n669) );
  XNOR2_X1 U727 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U728 ( .A(G107), .B(n671), .ZN(G9) );
  XNOR2_X1 U729 ( .A(G110), .B(n672), .ZN(G12) );
  XOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .Z(n675) );
  NAND2_X1 U731 ( .A1(n677), .A2(n673), .ZN(n674) );
  XNOR2_X1 U732 ( .A(n675), .B(n674), .ZN(G30) );
  NAND2_X1 U733 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n678), .B(KEYINPUT110), .ZN(n679) );
  XNOR2_X1 U735 ( .A(G146), .B(n679), .ZN(G48) );
  NOR2_X1 U736 ( .A1(n680), .A2(n682), .ZN(n681) );
  XOR2_X1 U737 ( .A(G113), .B(n681), .Z(G15) );
  NOR2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n685) );
  XNOR2_X1 U739 ( .A(G116), .B(KEYINPUT111), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n685), .B(n684), .ZN(G18) );
  XNOR2_X1 U741 ( .A(G125), .B(n686), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n687), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U743 ( .A(G134), .B(n688), .ZN(G36) );
  XOR2_X1 U744 ( .A(G140), .B(n689), .Z(G42) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  NAND2_X1 U746 ( .A1(n349), .A2(G469), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n706), .A2(n692), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n700), .A2(G475), .ZN(n696) );
  XOR2_X1 U749 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n693) );
  XNOR2_X1 U750 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U751 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n698) );
  NAND2_X1 U752 ( .A1(n349), .A2(G217), .ZN(n704) );
  INV_X1 U753 ( .A(KEYINPUT123), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U755 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U756 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U757 ( .A1(n708), .A2(G898), .ZN(n711) );
  NAND2_X1 U758 ( .A1(n709), .A2(n443), .ZN(n710) );
  NAND2_X1 U759 ( .A1(n711), .A2(n710), .ZN(n715) );
  OR2_X1 U760 ( .A1(n443), .A2(G898), .ZN(n713) );
  NAND2_X1 U761 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U762 ( .A(n715), .B(n714), .Z(G69) );
  XNOR2_X1 U763 ( .A(KEYINPUT84), .B(KEYINPUT124), .ZN(n718) );
  XNOR2_X1 U764 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U765 ( .A(n716), .B(n719), .ZN(n724) );
  INV_X1 U766 ( .A(n724), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U768 ( .A1(G953), .A2(n722), .ZN(n723) );
  XNOR2_X1 U769 ( .A(KEYINPUT125), .B(n723), .ZN(n728) );
  XNOR2_X1 U770 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n728), .A2(n727), .ZN(G72) );
  XNOR2_X1 U774 ( .A(n729), .B(G131), .ZN(G33) );
  XOR2_X1 U775 ( .A(G143), .B(n730), .Z(G45) );
  XNOR2_X1 U776 ( .A(n731), .B(G122), .ZN(G24) );
  XNOR2_X1 U777 ( .A(G119), .B(n732), .ZN(G21) );
  XNOR2_X1 U778 ( .A(G137), .B(KEYINPUT126), .ZN(n734) );
  XNOR2_X1 U779 ( .A(n734), .B(n733), .ZN(G39) );
endmodule

