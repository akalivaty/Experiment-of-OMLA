

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599;

  XNOR2_X1 U323 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n347) );
  NOR2_X1 U324 ( .A1(n586), .A2(n477), .ZN(n478) );
  NOR2_X1 U325 ( .A1(n546), .A2(n520), .ZN(n465) );
  XOR2_X1 U326 ( .A(n327), .B(n343), .Z(n552) );
  NOR2_X1 U327 ( .A1(n499), .A2(n504), .ZN(n345) );
  XNOR2_X1 U328 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n468) );
  XNOR2_X1 U329 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U330 ( .A(KEYINPUT99), .ZN(n353) );
  INV_X1 U331 ( .A(n386), .ZN(n387) );
  XNOR2_X1 U332 ( .A(n354), .B(n353), .ZN(n371) );
  XNOR2_X1 U333 ( .A(n307), .B(G120GAT), .ZN(n431) );
  XNOR2_X1 U334 ( .A(n388), .B(n387), .ZN(n389) );
  NAND2_X1 U335 ( .A1(n371), .A2(n373), .ZN(n372) );
  XNOR2_X1 U336 ( .A(n390), .B(n389), .ZN(n394) );
  XNOR2_X1 U337 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U338 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U339 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U340 ( .A(n322), .B(n321), .ZN(n327) );
  NOR2_X1 U341 ( .A1(n500), .A2(n499), .ZN(n587) );
  XOR2_X1 U342 ( .A(KEYINPUT92), .B(n373), .Z(n547) );
  INV_X1 U343 ( .A(n552), .ZN(n499) );
  XNOR2_X1 U344 ( .A(n501), .B(G176GAT), .ZN(n502) );
  XNOR2_X1 U345 ( .A(n490), .B(G134GAT), .ZN(n491) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n466) );
  XNOR2_X1 U347 ( .A(n503), .B(n502), .ZN(G1349GAT) );
  XNOR2_X1 U348 ( .A(n467), .B(n466), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G148GAT), .B(KEYINPUT88), .Z(n293) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G218GAT), .Z(n386) );
  XNOR2_X1 U351 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n291) );
  XNOR2_X1 U352 ( .A(n291), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U353 ( .A(n386), .B(n332), .ZN(n292) );
  XNOR2_X1 U354 ( .A(n293), .B(n292), .ZN(n298) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U356 ( .A(n294), .B(G204GAT), .ZN(n430) );
  XOR2_X1 U357 ( .A(n430), .B(KEYINPUT87), .Z(n296) );
  NAND2_X1 U358 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U359 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U360 ( .A(n298), .B(n297), .Z(n306) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(G162GAT), .Z(n300) );
  XNOR2_X1 U362 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n299) );
  XNOR2_X1 U363 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U364 ( .A(G141GAT), .B(n301), .Z(n368) );
  XOR2_X1 U365 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n303) );
  XNOR2_X1 U366 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n302) );
  XNOR2_X1 U367 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n368), .B(n304), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n496) );
  XOR2_X1 U370 ( .A(G43GAT), .B(G134GAT), .Z(n385) );
  XNOR2_X1 U371 ( .A(G99GAT), .B(G71GAT), .ZN(n307) );
  XNOR2_X1 U372 ( .A(n385), .B(n431), .ZN(n311) );
  INV_X1 U373 ( .A(n311), .ZN(n309) );
  AND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n310) );
  INV_X1 U375 ( .A(n310), .ZN(n308) );
  NAND2_X1 U376 ( .A1(n309), .A2(n308), .ZN(n313) );
  NAND2_X1 U377 ( .A1(n311), .A2(n310), .ZN(n312) );
  NAND2_X1 U378 ( .A1(n313), .A2(n312), .ZN(n315) );
  INV_X1 U379 ( .A(KEYINPUT20), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n322) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U382 ( .A(n316), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U383 ( .A(n360), .B(KEYINPUT83), .ZN(n320) );
  XOR2_X1 U384 ( .A(G176GAT), .B(KEYINPUT85), .Z(n318) );
  XNOR2_X1 U385 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n317) );
  XNOR2_X1 U386 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n324) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U390 ( .A(G190GAT), .B(KEYINPUT18), .Z(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n343) );
  XOR2_X1 U392 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n329) );
  XNOR2_X1 U393 ( .A(G204GAT), .B(KEYINPUT94), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n342) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G64GAT), .Z(n438) );
  INV_X1 U396 ( .A(n438), .ZN(n331) );
  INV_X1 U397 ( .A(n332), .ZN(n330) );
  NAND2_X1 U398 ( .A1(n331), .A2(n330), .ZN(n334) );
  NAND2_X1 U399 ( .A1(n438), .A2(n332), .ZN(n333) );
  NAND2_X1 U400 ( .A1(n334), .A2(n333), .ZN(n336) );
  AND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n338) );
  INV_X1 U403 ( .A(G92GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U405 ( .A(G36GAT), .B(G8GAT), .Z(n458) );
  XNOR2_X1 U406 ( .A(n458), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n504) );
  XOR2_X1 U410 ( .A(KEYINPUT97), .B(n345), .Z(n346) );
  NOR2_X1 U411 ( .A1(n496), .A2(n346), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n350) );
  NAND2_X1 U414 ( .A1(n496), .A2(n499), .ZN(n349) );
  XOR2_X1 U415 ( .A(n350), .B(n349), .Z(n508) );
  INV_X1 U416 ( .A(n508), .ZN(n566) );
  INV_X1 U417 ( .A(n504), .ZN(n549) );
  XNOR2_X1 U418 ( .A(KEYINPUT27), .B(n549), .ZN(n374) );
  NAND2_X1 U419 ( .A1(n566), .A2(n374), .ZN(n351) );
  NAND2_X1 U420 ( .A1(n352), .A2(n351), .ZN(n354) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n356) );
  XNOR2_X1 U422 ( .A(G120GAT), .B(KEYINPUT91), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U424 ( .A(n357), .B(G85GAT), .Z(n359) );
  XOR2_X1 U425 ( .A(G148GAT), .B(G57GAT), .Z(n439) );
  XNOR2_X1 U426 ( .A(G134GAT), .B(n439), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n364) );
  XOR2_X1 U428 ( .A(G29GAT), .B(G1GAT), .Z(n452) );
  XOR2_X1 U429 ( .A(n360), .B(n452), .Z(n362) );
  NAND2_X1 U430 ( .A1(G225GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U432 ( .A(n364), .B(n363), .Z(n370) );
  XOR2_X1 U433 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n366) );
  XNOR2_X1 U434 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n372), .B(KEYINPUT100), .ZN(n378) );
  NAND2_X1 U439 ( .A1(n547), .A2(n374), .ZN(n482) );
  XOR2_X1 U440 ( .A(KEYINPUT86), .B(n499), .Z(n375) );
  NOR2_X1 U441 ( .A1(n482), .A2(n375), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n496), .B(KEYINPUT28), .ZN(n554) );
  INV_X1 U443 ( .A(n554), .ZN(n533) );
  NAND2_X1 U444 ( .A1(n376), .A2(n533), .ZN(n377) );
  NAND2_X1 U445 ( .A1(n378), .A2(n377), .ZN(n518) );
  XOR2_X1 U446 ( .A(G106GAT), .B(G162GAT), .Z(n380) );
  XNOR2_X1 U447 ( .A(G190GAT), .B(G99GAT), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U449 ( .A(G85GAT), .B(G92GAT), .Z(n443) );
  XNOR2_X1 U450 ( .A(n381), .B(n443), .ZN(n383) );
  XOR2_X1 U451 ( .A(G29GAT), .B(G36GAT), .Z(n382) );
  XNOR2_X1 U452 ( .A(n383), .B(n382), .ZN(n390) );
  XNOR2_X1 U453 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n384), .B(KEYINPUT69), .ZN(n447) );
  XNOR2_X1 U455 ( .A(n447), .B(n385), .ZN(n388) );
  XOR2_X1 U456 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n392) );
  NAND2_X1 U457 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  XOR2_X1 U458 ( .A(n392), .B(n391), .Z(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U460 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n396) );
  XNOR2_X1 U461 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n397), .B(KEYINPUT72), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n400) );
  NAND2_X1 U465 ( .A1(n400), .A2(KEYINPUT102), .ZN(n403) );
  INV_X1 U466 ( .A(n400), .ZN(n474) );
  INV_X1 U467 ( .A(KEYINPUT102), .ZN(n401) );
  NAND2_X1 U468 ( .A1(n474), .A2(n401), .ZN(n402) );
  NAND2_X1 U469 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n404), .B(KEYINPUT36), .ZN(n596) );
  XOR2_X1 U471 ( .A(KEYINPUT80), .B(KEYINPUT76), .Z(n406) );
  XNOR2_X1 U472 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n414) );
  NAND2_X1 U474 ( .A1(G231GAT), .A2(G233GAT), .ZN(n412) );
  XOR2_X1 U475 ( .A(G211GAT), .B(G78GAT), .Z(n408) );
  XNOR2_X1 U476 ( .A(G71GAT), .B(G155GAT), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U478 ( .A(G183GAT), .B(G127GAT), .Z(n409) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n426) );
  XOR2_X1 U482 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n416) );
  XNOR2_X1 U483 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U485 ( .A(KEYINPUT13), .B(G64GAT), .Z(n418) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(G57GAT), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n424) );
  XNOR2_X1 U489 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n422) );
  XNOR2_X1 U490 ( .A(G15GAT), .B(G22GAT), .ZN(n421) );
  XOR2_X1 U491 ( .A(n421), .B(KEYINPUT70), .Z(n451) );
  XNOR2_X1 U492 ( .A(n422), .B(n451), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U494 ( .A(n426), .B(n425), .Z(n515) );
  AND2_X1 U495 ( .A1(n596), .A2(n515), .ZN(n427) );
  AND2_X1 U496 ( .A1(n518), .A2(n427), .ZN(n429) );
  XOR2_X1 U497 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n428) );
  XNOR2_X1 U498 ( .A(n429), .B(n428), .ZN(n546) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n436) );
  XOR2_X1 U500 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n433) );
  NAND2_X1 U501 ( .A1(G230GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U502 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U503 ( .A(n434), .B(KEYINPUT13), .Z(n435) );
  XNOR2_X1 U504 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U505 ( .A(n437), .B(KEYINPUT31), .Z(n442) );
  XNOR2_X1 U506 ( .A(n438), .B(KEYINPUT71), .ZN(n440) );
  XOR2_X1 U507 ( .A(n444), .B(n443), .Z(n590) );
  XOR2_X1 U508 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n450) );
  XOR2_X1 U509 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n446) );
  XNOR2_X1 U510 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n452), .B(n451), .ZN(n454) );
  NAND2_X1 U515 ( .A1(G229GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n462) );
  XOR2_X1 U517 ( .A(G141GAT), .B(G197GAT), .Z(n456) );
  XNOR2_X1 U518 ( .A(G43GAT), .B(G50GAT), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U520 ( .A(n457), .B(G113GAT), .Z(n460) );
  XNOR2_X1 U521 ( .A(G169GAT), .B(n458), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U523 ( .A(n462), .B(n461), .Z(n463) );
  XOR2_X1 U524 ( .A(n464), .B(n463), .Z(n568) );
  OR2_X1 U525 ( .A1(n590), .A2(n568), .ZN(n520) );
  XOR2_X1 U526 ( .A(KEYINPUT38), .B(n465), .Z(n532) );
  OR2_X1 U527 ( .A1(n532), .A2(n499), .ZN(n467) );
  INV_X1 U528 ( .A(n515), .ZN(n593) );
  NAND2_X1 U529 ( .A1(n596), .A2(n593), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n590), .A2(n470), .ZN(n471) );
  XNOR2_X1 U531 ( .A(KEYINPUT112), .B(n471), .ZN(n472) );
  AND2_X1 U532 ( .A1(n568), .A2(n472), .ZN(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT113), .B(n473), .ZN(n480) );
  INV_X1 U534 ( .A(n474), .ZN(n586) );
  INV_X1 U535 ( .A(n568), .ZN(n580) );
  XOR2_X1 U536 ( .A(KEYINPUT41), .B(n590), .Z(n571) );
  NAND2_X1 U537 ( .A1(n580), .A2(n571), .ZN(n475) );
  XNOR2_X1 U538 ( .A(KEYINPUT46), .B(n475), .ZN(n476) );
  NAND2_X1 U539 ( .A1(n476), .A2(n515), .ZN(n477) );
  XNOR2_X1 U540 ( .A(KEYINPUT47), .B(n478), .ZN(n479) );
  AND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT48), .B(n481), .ZN(n493) );
  NOR2_X1 U543 ( .A1(n493), .A2(n482), .ZN(n567) );
  AND2_X1 U544 ( .A1(n567), .A2(n552), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(KEYINPUT114), .ZN(n484) );
  NAND2_X1 U546 ( .A1(n484), .A2(n533), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n485), .B(KEYINPUT115), .ZN(n563) );
  NAND2_X1 U548 ( .A1(n563), .A2(n593), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n487) );
  XNOR2_X1 U550 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1342GAT) );
  NAND2_X1 U553 ( .A1(n563), .A2(n586), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n490) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1343GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT106), .B(n571), .ZN(n562) );
  XOR2_X1 U557 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n498) );
  NOR2_X1 U558 ( .A1(n493), .A2(n504), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n494), .B(KEYINPUT54), .ZN(n495) );
  INV_X1 U560 ( .A(n547), .ZN(n529) );
  NAND2_X1 U561 ( .A1(n495), .A2(n529), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n509), .A2(n496), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n500) );
  NAND2_X1 U564 ( .A1(n562), .A2(n587), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n501) );
  NOR2_X1 U566 ( .A1(n532), .A2(n504), .ZN(n507) );
  INV_X1 U567 ( .A(G36GAT), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n511) );
  NOR2_X1 U571 ( .A1(n509), .A2(n508), .ZN(n597) );
  NAND2_X1 U572 ( .A1(n597), .A2(n580), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n512), .B(KEYINPUT59), .ZN(n514) );
  XOR2_X1 U575 ( .A(G197GAT), .B(KEYINPUT125), .Z(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1352GAT) );
  NOR2_X1 U577 ( .A1(n586), .A2(n515), .ZN(n517) );
  XNOR2_X1 U578 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(n519) );
  NAND2_X1 U580 ( .A1(n519), .A2(n518), .ZN(n535) );
  NOR2_X1 U581 ( .A1(n520), .A2(n535), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n527), .A2(n547), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n521), .B(KEYINPUT34), .ZN(n522) );
  XNOR2_X1 U584 ( .A(G1GAT), .B(n522), .ZN(G1324GAT) );
  NAND2_X1 U585 ( .A1(n527), .A2(n549), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n525) );
  NAND2_X1 U588 ( .A1(n527), .A2(n552), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U590 ( .A(G15GAT), .B(n526), .Z(G1326GAT) );
  NAND2_X1 U591 ( .A1(n554), .A2(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U593 ( .A1(n532), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1328GAT) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(G50GAT), .B(n534), .Z(G1331GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n537) );
  NAND2_X1 U599 ( .A1(n568), .A2(n562), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n545), .A2(n535), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n542), .A2(n547), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G57GAT), .B(n538), .ZN(G1332GAT) );
  XOR2_X1 U604 ( .A(G64GAT), .B(KEYINPUT107), .Z(n540) );
  NAND2_X1 U605 ( .A1(n542), .A2(n549), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1333GAT) );
  NAND2_X1 U607 ( .A1(n542), .A2(n552), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n541), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U609 ( .A(G78GAT), .B(KEYINPUT43), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n554), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1335GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n547), .A2(n555), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G85GAT), .B(n548), .ZN(G1336GAT) );
  XNOR2_X1 U615 ( .A(G92GAT), .B(KEYINPUT108), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n555), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1337GAT) );
  NAND2_X1 U618 ( .A1(n555), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n557) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(n558), .B(KEYINPUT110), .Z(n560) );
  XNOR2_X1 U624 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1339GAT) );
  NAND2_X1 U626 ( .A1(n580), .A2(n563), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U628 ( .A(G120GAT), .B(KEYINPUT49), .Z(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1341GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n570) );
  NOR2_X1 U632 ( .A1(n568), .A2(n570), .ZN(n569) );
  XOR2_X1 U633 ( .A(G141GAT), .B(n569), .Z(G1344GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n573) );
  INV_X1 U635 ( .A(n570), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G148GAT), .B(n574), .ZN(G1345GAT) );
  XOR2_X1 U639 ( .A(G155GAT), .B(KEYINPUT119), .Z(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n593), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1346GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n586), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT120), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G162GAT), .B(n579), .ZN(G1347GAT) );
  XNOR2_X1 U645 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n587), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1348GAT) );
  NAND2_X1 U648 ( .A1(n587), .A2(n593), .ZN(n584) );
  XOR2_X1 U649 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT58), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G190GAT), .B(n589), .ZN(G1351GAT) );
  XOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT61), .Z(n592) );
  NAND2_X1 U656 ( .A1(n597), .A2(n590), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1353GAT) );
  XOR2_X1 U658 ( .A(G211GAT), .B(KEYINPUT127), .Z(n595) );
  NAND2_X1 U659 ( .A1(n597), .A2(n593), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n595), .B(n594), .ZN(G1354GAT) );
  NAND2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U662 ( .A(n598), .B(KEYINPUT62), .ZN(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

