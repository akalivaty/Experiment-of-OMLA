//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G101), .A3(new_n465), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT3), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n481), .A2(G137), .A3(new_n465), .A4(new_n468), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n465), .A3(new_n468), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n465), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n481), .A2(G2105), .A3(new_n468), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n495), .B2(G124), .ZN(new_n496));
  XOR2_X1   g071(.A(new_n496), .B(KEYINPUT70), .Z(G162));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AND4_X1   g074(.A1(new_n465), .A2(new_n499), .A3(new_n468), .A4(new_n470), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n481), .A2(G138), .A3(new_n465), .A4(new_n468), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n481), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n502), .A2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n512), .A2(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT72), .B(G89), .Z(new_n531));
  OAI211_X1 g106(.A(new_n529), .B(new_n530), .C1(new_n510), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(G168));
  AND2_X1   g108(.A1(new_n526), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n535), .A2(new_n516), .B1(new_n510), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  XNOR2_X1  g113(.A(KEYINPUT73), .B(G43), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n526), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n508), .A2(new_n509), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(KEYINPUT5), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(G81), .A2(new_n541), .B1(new_n547), .B2(G651), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n512), .B2(new_n557), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  OAI211_X1 g136(.A(KEYINPUT75), .B(new_n561), .C1(new_n512), .C2(new_n557), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n545), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(G91), .A2(new_n541), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n541), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n523), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n508), .A2(new_n509), .A3(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n508), .A2(new_n509), .A3(new_n578), .A4(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n545), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n516), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT77), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT78), .B(G47), .Z(new_n589));
  AOI22_X1  g164(.A1(new_n526), .A2(new_n589), .B1(G85), .B2(new_n541), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(G290));
  AND3_X1   g166(.A1(new_n508), .A2(new_n509), .A3(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n526), .A2(G54), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n516), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G321));
  NOR2_X1   g176(.A1(G286), .A2(new_n598), .ZN(new_n602));
  XNOR2_X1  g177(.A(G299), .B(KEYINPUT79), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n598), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n598), .ZN(G280));
  AND3_X1   g180(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g187(.A1(new_n479), .A2(new_n463), .A3(new_n465), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2100), .Z(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT81), .B(G2096), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n465), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n485), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n493), .A2(new_n494), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n622), .A2(KEYINPUT80), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT80), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n616), .B1(new_n617), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n617), .B2(new_n626), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT82), .Z(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n638), .B(new_n640), .Z(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G14), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n641), .B2(new_n643), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(KEYINPUT17), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n653), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n654), .B(KEYINPUT86), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n656), .B(new_n660), .C1(new_n658), .C2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT87), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G33), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G139), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n485), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT94), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  OAI22_X1  g269(.A1(new_n692), .A2(new_n693), .B1(new_n465), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT95), .Z(new_n696));
  OAI21_X1  g271(.A(new_n685), .B1(new_n696), .B2(new_n684), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT96), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n698), .A2(G2072), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT100), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT99), .B(KEYINPUT26), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n486), .A2(G141), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n479), .A2(G105), .A3(new_n465), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n495), .A2(G129), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(KEYINPUT98), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(KEYINPUT98), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n684), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n684), .B2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G2084), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n684), .B1(KEYINPUT24), .B2(G34), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(KEYINPUT24), .B2(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n483), .B2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n716), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G2072), .B2(new_n698), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n701), .A2(KEYINPUT101), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(KEYINPUT101), .B1(new_n701), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G23), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n574), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n725), .A2(G6), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G305), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT32), .B(G1981), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G22), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G166), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1971), .Z(new_n740));
  OAI211_X1 g315(.A(new_n734), .B(new_n740), .C1(new_n731), .C2(new_n733), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT34), .ZN(new_n742));
  MUX2_X1   g317(.A(G24), .B(G290), .S(new_n737), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1986), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n684), .A2(G25), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT88), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n495), .A2(G119), .ZN(new_n747));
  NOR2_X1   g322(.A1(G95), .A2(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT89), .Z(new_n749));
  INV_X1    g324(.A(G107), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n469), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n486), .A2(G131), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n744), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n741), .A2(KEYINPUT34), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n742), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT36), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n725), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n725), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT102), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1966), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n684), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n725), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n725), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(new_n770), .B2(G1961), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G1961), .B2(new_n770), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n737), .A2(G19), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n549), .B2(new_n737), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1341), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n717), .B2(new_n720), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT92), .Z(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n597), .B2(new_n725), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G29), .B2(new_n626), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n764), .A2(new_n772), .A3(new_n776), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n735), .A2(G20), .A3(new_n736), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(G299), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n725), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n684), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n684), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n793), .C1(new_n714), .C2(new_n715), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n684), .A2(G26), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n495), .A2(G128), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n465), .A2(G116), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n486), .A2(G140), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT93), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n783), .A2(new_n794), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G35), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G162), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT29), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G2090), .Z(new_n810));
  NAND3_X1  g385(.A1(new_n760), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n723), .A2(new_n724), .A3(new_n811), .ZN(G311));
  INV_X1    g387(.A(new_n724), .ZN(new_n813));
  INV_X1    g388(.A(new_n811), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n701), .A2(KEYINPUT101), .A3(new_n722), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(G150));
  NAND2_X1  g391(.A1(new_n606), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n526), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(new_n516), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT103), .B(G93), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n541), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n549), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n540), .A2(new_n548), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n818), .B(new_n829), .Z(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n831), .A2(new_n832), .A3(G860), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n826), .A2(G860), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(new_n835), .ZN(G145));
  NAND2_X1  g411(.A1(new_n710), .A2(new_n711), .ZN(new_n837));
  INV_X1    g412(.A(new_n708), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n695), .B(KEYINPUT95), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n696), .A2(new_n712), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n844));
  INV_X1    g419(.A(new_n500), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n847));
  INV_X1    g422(.A(new_n506), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT104), .B1(new_n502), .B2(new_n506), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n802), .B(new_n851), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n841), .A3(new_n842), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n495), .A2(G130), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n465), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n486), .A2(G142), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n753), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n753), .A2(new_n863), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n865), .A2(new_n866), .A3(new_n614), .ZN(new_n867));
  INV_X1    g442(.A(new_n614), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n747), .A2(new_n752), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT105), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n862), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n614), .B1(new_n865), .B2(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n868), .A3(new_n864), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n873), .A2(new_n857), .A3(new_n861), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT106), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n856), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n877), .A2(new_n876), .B1(new_n853), .B2(new_n855), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G162), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n626), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n880), .B2(new_n881), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n881), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n878), .A2(new_n879), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n884), .B(new_n889), .C1(new_n890), .C2(new_n856), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  AND4_X1   g467(.A1(KEYINPUT40), .A2(new_n891), .A3(new_n892), .A4(new_n887), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n888), .A2(new_n893), .ZN(G395));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n824), .B2(G868), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT107), .B1(new_n606), .B2(G299), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n786), .A2(new_n597), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n606), .A2(G299), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n897), .A2(new_n899), .A3(KEYINPUT41), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n829), .B(new_n609), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT42), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(KEYINPUT42), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G166), .B(KEYINPUT108), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(G305), .ZN(new_n914));
  XNOR2_X1  g489(.A(G290), .B(new_n574), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n598), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n910), .A2(new_n911), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n896), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n917), .A2(new_n919), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(KEYINPUT109), .B2(new_n921), .ZN(G295));
  AOI21_X1  g497(.A(new_n920), .B1(KEYINPUT109), .B2(new_n921), .ZN(G331));
  AOI21_X1  g498(.A(G301), .B1(new_n825), .B2(new_n828), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n825), .A2(G301), .A3(new_n828), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(G168), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G286), .B1(new_n928), .B2(new_n924), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n901), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n905), .A2(new_n927), .A3(new_n929), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n916), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n892), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n916), .B1(new_n931), .B2(new_n932), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n934), .A2(KEYINPUT43), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n927), .B(new_n929), .C1(KEYINPUT110), .C2(new_n904), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n903), .A2(KEYINPUT110), .A3(new_n904), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n934), .B1(new_n918), .B2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n936), .B(KEYINPUT44), .C1(new_n937), .C2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n934), .B2(new_n935), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n918), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n945), .A2(new_n937), .A3(new_n892), .A4(new_n933), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g524(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n944), .C2(new_n946), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(G397));
  AND3_X1   g526(.A1(new_n482), .A2(new_n480), .A3(G40), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n475), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n502), .B2(new_n506), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n953), .A2(new_n955), .A3(G2067), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n957));
  INV_X1    g532(.A(new_n953), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n959), .B(new_n954), .C1(new_n502), .C2(new_n506), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n961), .B2(new_n780), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(new_n597), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n788), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n953), .B1(new_n965), .B2(new_n955), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT45), .A4(new_n954), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT56), .B(G2072), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G299), .A2(KEYINPUT57), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT57), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n560), .A2(new_n971), .A3(new_n562), .A4(new_n566), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n964), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n963), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n964), .A2(new_n969), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n966), .A2(new_n967), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT58), .B(G1341), .Z(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n953), .B2(new_n955), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT118), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n981), .C1(new_n953), .C2(new_n955), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n986), .A2(KEYINPUT59), .A3(new_n549), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT59), .B1(new_n986), .B2(new_n549), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n977), .A2(new_n973), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT61), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n961), .A2(new_n780), .ZN(new_n993));
  INV_X1    g568(.A(new_n956), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(KEYINPUT60), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n606), .B1(new_n962), .B2(KEYINPUT60), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n962), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n989), .B(new_n992), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT119), .B1(new_n990), .B2(new_n991), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n977), .A2(new_n1004), .A3(KEYINPUT61), .A4(new_n973), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n978), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n583), .A2(G651), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n523), .A2(G48), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n576), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G1981), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n580), .A2(new_n584), .A3(new_n1012), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1011), .A2(new_n1013), .A3(KEYINPUT49), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT49), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n955), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n958), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n574), .A2(G1976), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1017), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1020), .B(new_n1021), .C1(new_n955), .C2(new_n953), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1016), .A2(new_n1019), .B1(KEYINPUT52), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n574), .A2(G1976), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1022), .A2(KEYINPUT52), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n961), .A2(G2090), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1971), .B1(new_n966), .B2(new_n967), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1021), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(G166), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT55), .B(G8), .C1(new_n514), .C2(new_n517), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1033), .A2(KEYINPUT114), .A3(new_n1034), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(G8), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1027), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n955), .A2(new_n965), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT45), .B(new_n954), .C1(new_n502), .C2(new_n506), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n958), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT117), .B(G2084), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n957), .A2(new_n958), .A3(new_n960), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1032), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G168), .A2(new_n1017), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1041), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1966), .B1(new_n966), .B2(new_n1043), .ZN(new_n1052));
  AND4_X1   g627(.A1(new_n958), .A2(new_n957), .A3(new_n960), .A4(new_n1047), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT122), .B(new_n1021), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1017), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(KEYINPUT122), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1051), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1040), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n966), .A2(new_n967), .A3(new_n792), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n965), .B1(new_n851), .B2(G1384), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n473), .B2(G2105), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n952), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n967), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n961), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1064), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G171), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1062), .A2(new_n1063), .B1(new_n1070), .B2(new_n961), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n966), .A2(KEYINPUT53), .A3(new_n792), .A4(new_n1043), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(G301), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(KEYINPUT54), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT125), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1073), .A2(new_n1079), .A3(KEYINPUT54), .A4(new_n1076), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT124), .B1(new_n1072), .B2(G171), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1074), .A2(new_n1084), .A3(G301), .A4(new_n1069), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1078), .A2(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1007), .A2(new_n1061), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(G288), .A2(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1013), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1019), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n966), .A2(new_n967), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1098), .A2(G1971), .B1(G2090), .B2(new_n961), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1099), .B2(G8), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1057), .A2(new_n1023), .A3(G168), .A4(new_n1025), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT63), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1039), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1057), .A2(new_n1104), .A3(G168), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1105), .B2(new_n1035), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1096), .B(new_n1102), .C1(new_n1106), .C2(new_n1026), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1027), .A2(new_n1035), .A3(new_n1108), .A4(new_n1039), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1059), .A2(new_n1112), .A3(new_n1060), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1089), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n869), .B(new_n755), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n802), .A2(G2067), .ZN(new_n1118));
  INV_X1    g693(.A(G2067), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n797), .A2(new_n1119), .A3(new_n801), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1118), .A2(KEYINPUT112), .A3(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n712), .B(G1996), .ZN(new_n1126));
  XOR2_X1   g701(.A(G290), .B(G1986), .Z(new_n1127));
  NAND4_X1  g702(.A1(new_n1117), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1065), .A2(new_n953), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1115), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n839), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1129), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1133), .A2(new_n1134), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1129), .A2(new_n979), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT46), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1136), .B(new_n1139), .Z(new_n1140));
  OR3_X1    g715(.A1(new_n1135), .A2(new_n1140), .A3(KEYINPUT47), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT47), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1126), .A2(new_n1125), .A3(new_n755), .A4(new_n869), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1134), .B1(new_n1144), .B2(new_n1120), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1117), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1129), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1134), .A2(G1986), .A3(G290), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT48), .Z(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1143), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1131), .A2(new_n1132), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1130), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1089), .B2(new_n1114), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT127), .B1(new_n1155), .B2(new_n1151), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g732(.A1(new_n885), .A2(new_n887), .ZN(new_n1159));
  INV_X1    g733(.A(G319), .ZN(new_n1160));
  NOR2_X1   g734(.A1(G227), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n682), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n1162), .B1(new_n646), .B2(new_n648), .ZN(new_n1163));
  AND3_X1   g737(.A1(new_n1159), .A2(new_n1163), .A3(new_n947), .ZN(G308));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1163), .A3(new_n947), .ZN(G225));
endmodule


