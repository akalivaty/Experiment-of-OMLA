//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT64), .B1(new_n203), .B2(G146), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n200), .B(new_n202), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G143), .B2(new_n199), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n210), .B2(new_n201), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n215));
  XNOR2_X1  g029(.A(G104), .B(G107), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G107), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT76), .A3(G101), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n219), .A3(G104), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n225), .A2(new_n227), .A3(new_n222), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n218), .A2(new_n224), .B1(new_n228), .B2(new_n217), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n206), .A2(new_n211), .A3(KEYINPUT67), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n214), .A2(new_n229), .A3(KEYINPUT10), .A4(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(new_n227), .A3(new_n222), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n225), .A2(new_n227), .A3(new_n217), .A4(new_n222), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n199), .B2(G143), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n237), .A2(new_n238), .B1(G143), .B2(new_n199), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n242), .A2(new_n240), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n239), .A2(new_n241), .B1(new_n243), .B2(new_n208), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n232), .A2(new_n245), .A3(G101), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n235), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n250));
  INV_X1    g064(.A(new_n206), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n237), .A2(new_n238), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n252), .A2(new_n200), .B1(G128), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT76), .B1(new_n223), .B2(G101), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n215), .B(new_n217), .C1(new_n220), .C2(new_n222), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n234), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT77), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n210), .A2(new_n201), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n206), .B1(new_n239), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n229), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT10), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(KEYINPUT78), .B(KEYINPUT10), .C1(new_n259), .C2(new_n263), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n198), .B(new_n249), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n218), .A2(new_n224), .ZN(new_n269));
  AND4_X1   g083(.A1(new_n260), .A2(new_n262), .A3(new_n234), .A4(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n260), .B1(new_n229), .B2(new_n262), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n229), .A2(new_n212), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT12), .B(new_n197), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n259), .B2(new_n263), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n198), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT68), .B(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G227), .ZN(new_n281));
  XOR2_X1   g095(.A(G110), .B(G140), .Z(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n249), .B1(new_n266), .B2(new_n267), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n197), .ZN(new_n286));
  INV_X1    g100(.A(new_n283), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n268), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT79), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT78), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n264), .A2(new_n250), .A3(new_n265), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n248), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n283), .B1(new_n296), .B2(new_n198), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n286), .A2(new_n297), .B1(new_n279), .B2(new_n283), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n292), .B(G469), .C1(new_n298), .C2(G902), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT80), .B(G469), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n287), .B1(new_n286), .B2(new_n268), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n268), .A2(new_n278), .A3(new_n287), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n291), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  OAI21_X1  g121(.A(G221), .B1(new_n307), .B2(G902), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT2), .B(G113), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G119), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT66), .A3(G116), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(G119), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n314), .A2(new_n317), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT5), .A4(new_n320), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n316), .A2(KEYINPUT5), .A3(G119), .ZN(new_n323));
  INV_X1    g137(.A(G113), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n269), .A2(new_n321), .A3(new_n234), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n235), .A2(new_n246), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n329), .A2(new_n330), .A3(new_n313), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n313), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n327), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G122), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT81), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT6), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n206), .A2(new_n211), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n252), .A2(new_n241), .A3(new_n200), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n208), .A2(new_n240), .A3(new_n242), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G224), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT84), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n344), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n334), .A2(KEYINPUT82), .A3(new_n336), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n327), .B(new_n335), .C1(new_n328), .C2(new_n333), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT82), .B1(new_n334), .B2(new_n336), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n351), .A2(KEYINPUT6), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT83), .A4(new_n350), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n338), .B(new_n348), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n346), .A2(KEYINPUT86), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n340), .B2(new_n343), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT7), .B1(new_n345), .B2(G953), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n361), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n359), .B(new_n363), .C1(new_n340), .C2(new_n343), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n322), .A2(KEYINPUT85), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n325), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n322), .A2(KEYINPUT85), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n269), .A2(new_n234), .A3(new_n321), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n321), .A2(new_n326), .ZN(new_n371));
  OAI22_X1  g185(.A1(new_n369), .A2(new_n370), .B1(new_n371), .B2(new_n229), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n335), .B(KEYINPUT8), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n374), .A3(KEYINPUT87), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n351), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT87), .B1(new_n365), .B2(new_n374), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n300), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n312), .B1(new_n358), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n338), .ZN(new_n380));
  INV_X1    g194(.A(new_n348), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT83), .B1(new_n382), .B2(new_n355), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n352), .A2(new_n349), .A3(new_n353), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n380), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n378), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n311), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n310), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n221), .ZN(new_n390));
  INV_X1    g204(.A(G953), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT68), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  INV_X1    g208(.A(G237), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n392), .A2(new_n394), .A3(G214), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n203), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n280), .A2(G143), .A3(G214), .A4(new_n395), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT18), .A3(G131), .ZN(new_n400));
  INV_X1    g214(.A(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G125), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n339), .A2(G140), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n199), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(new_n398), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n397), .A2(new_n398), .A3(new_n195), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n195), .B1(new_n397), .B2(new_n398), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n399), .A2(KEYINPUT17), .A3(G131), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT16), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n339), .A2(KEYINPUT16), .A3(G140), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G146), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G146), .B1(new_n413), .B2(new_n414), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n390), .B(new_n408), .C1(new_n411), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n399), .A2(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n397), .A2(new_n398), .A3(new_n195), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n418), .B(new_n412), .C1(new_n425), .C2(KEYINPUT17), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(KEYINPUT88), .A3(new_n390), .A4(new_n408), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n404), .B(KEYINPUT19), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n416), .B1(new_n429), .B2(new_n199), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n390), .B1(new_n431), .B2(new_n408), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n435));
  NOR2_X1   g249(.A1(G475), .A2(G902), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT20), .A4(new_n436), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n435), .A2(KEYINPUT20), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(KEYINPUT20), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n432), .B1(new_n422), .B2(new_n427), .ZN(new_n440));
  INV_X1    g254(.A(new_n436), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n390), .B1(new_n426), .B2(new_n408), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n422), .B2(new_n427), .ZN(new_n444));
  OAI21_X1  g258(.A(G475), .B1(new_n444), .B2(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G952), .ZN(new_n447));
  AOI211_X1 g261(.A(G953), .B(new_n447), .C1(G234), .C2(G237), .ZN(new_n448));
  AOI211_X1 g262(.A(new_n300), .B(new_n280), .C1(G234), .C2(G237), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(G898), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n188), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n316), .A2(G122), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G116), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n456), .A3(new_n219), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n454), .B2(KEYINPUT14), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(G116), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT14), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n454), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n453), .B(new_n457), .C1(new_n219), .C2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n452), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n466), .A2(G128), .A3(new_n203), .A4(new_n467), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(G134), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n452), .A2(KEYINPUT91), .A3(new_n188), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n454), .A2(new_n456), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G107), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n457), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n188), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n471), .A2(new_n472), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n465), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n307), .A2(new_n481), .A3(G953), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT93), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n482), .B(KEYINPUT93), .Z(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n465), .A3(new_n479), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT94), .ZN(new_n487));
  OR3_X1    g301(.A1(new_n480), .A2(KEYINPUT94), .A3(new_n483), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n300), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT95), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT95), .A4(new_n300), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n489), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n446), .A2(new_n451), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n306), .A2(new_n308), .A3(new_n388), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n188), .A2(G137), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n190), .A2(G134), .ZN(new_n502));
  OAI21_X1  g316(.A(G131), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n196), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n214), .A2(new_n504), .A3(new_n230), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n244), .A2(new_n197), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n333), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n333), .A3(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n500), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT71), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n280), .A2(G210), .A3(new_n395), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(KEYINPUT29), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n506), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n504), .A2(new_n212), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n506), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n508), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n510), .ZN(new_n528));
  INV_X1    g342(.A(new_n520), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n508), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n505), .A2(KEYINPUT28), .A3(new_n333), .A4(new_n506), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n514), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n530), .B(new_n531), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n521), .A2(new_n300), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G472), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n522), .A2(new_n508), .A3(new_n526), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n520), .A2(new_n510), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT31), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n510), .A2(new_n500), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n533), .A2(new_n532), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n529), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n527), .A2(new_n520), .A3(new_n510), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT70), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n542), .A2(new_n545), .A3(new_n550), .A4(new_n547), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n539), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI211_X1 g368(.A(KEYINPUT32), .B(new_n539), .C1(new_n549), .C2(new_n551), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n537), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G234), .ZN(new_n557));
  OAI21_X1  g371(.A(G217), .B1(new_n557), .B2(G902), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT72), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n404), .A2(new_n199), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT73), .B1(new_n318), .B2(G128), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT73), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n201), .A3(G119), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n318), .A2(G128), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT24), .B(G110), .Z(new_n567));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n318), .B2(G128), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n570));
  INV_X1    g384(.A(G110), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(new_n565), .ZN(new_n572));
  OAI22_X1  g386(.A1(new_n566), .A2(new_n567), .B1(new_n572), .B2(KEYINPUT74), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n415), .B(new_n561), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n567), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n565), .A3(new_n570), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G110), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n576), .B(new_n578), .C1(new_n416), .C2(new_n417), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n579), .A3(new_n583), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n560), .B1(new_n587), .B2(G902), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n559), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n558), .A2(new_n300), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT75), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n556), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n499), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(new_n217), .ZN(G3));
  AOI21_X1  g412(.A(G902), .B1(new_n549), .B2(new_n551), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n552), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n306), .A2(new_n602), .A3(new_n595), .A4(new_n308), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n486), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n483), .B2(new_n480), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n486), .A2(new_n605), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT33), .B1(new_n487), .B2(new_n488), .ZN(new_n610));
  OAI211_X1 g424(.A(G478), .B(new_n300), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n446), .ZN(new_n614));
  INV_X1    g428(.A(new_n451), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n358), .A2(new_n378), .A3(new_n312), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n311), .B1(new_n385), .B2(new_n386), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n309), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n603), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n445), .B(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n437), .A2(new_n442), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n497), .ZN(new_n625));
  OR3_X1    g439(.A1(new_n618), .A2(new_n625), .A3(KEYINPUT98), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT98), .B1(new_n618), .B2(new_n625), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n603), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NOR2_X1   g444(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n580), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n591), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n590), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n602), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n499), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NAND2_X1  g454(.A1(new_n549), .A2(new_n551), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n538), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT32), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n552), .A2(new_n553), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n635), .B1(new_n645), .B2(new_n537), .ZN(new_n646));
  INV_X1    g460(.A(new_n308), .ZN(new_n647));
  OAI21_X1  g461(.A(G469), .B1(new_n298), .B2(G902), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n294), .A2(new_n295), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n198), .B1(new_n649), .B2(new_n249), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n197), .B(new_n248), .C1(new_n294), .C2(new_n295), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n283), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n268), .A2(new_n278), .A3(new_n287), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n648), .A2(KEYINPUT79), .B1(new_n654), .B2(new_n302), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n647), .B1(new_n655), .B2(new_n299), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n448), .B1(new_n449), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n625), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n646), .A2(new_n656), .A3(new_n388), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n658), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n528), .A2(new_n520), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n509), .A2(new_n510), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n300), .B1(new_n667), .B2(new_n520), .ZN(new_n668));
  OAI21_X1  g482(.A(G472), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n645), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n379), .A2(new_n387), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n446), .A2(new_n497), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n635), .A2(new_n309), .ZN(new_n676));
  NOR4_X1   g490(.A1(new_n671), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n664), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  INV_X1    g494(.A(new_n658), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n613), .A2(new_n446), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n646), .A2(new_n656), .A3(new_n388), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT99), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n306), .A2(new_n308), .A3(new_n388), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n556), .A2(new_n636), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n683), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT100), .B(G146), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G48));
  NOR2_X1   g507(.A1(new_n618), .A2(new_n614), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n305), .B(new_n308), .C1(new_n654), .C2(new_n290), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n694), .A2(new_n556), .A3(new_n595), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND3_X1  g513(.A1(new_n556), .A2(new_n696), .A3(new_n595), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n626), .B2(new_n627), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n316), .ZN(G18));
  OAI21_X1  g516(.A(new_n309), .B1(new_n616), .B2(new_n617), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n556), .A3(new_n498), .A4(new_n636), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  OAI211_X1 g520(.A(new_n513), .B(new_n529), .C1(new_n511), .C2(new_n515), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n542), .A3(new_n547), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n538), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n709), .B(new_n593), .C1(new_n599), .C2(new_n600), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n446), .A2(new_n711), .A3(new_n497), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n711), .B1(new_n446), .B2(new_n497), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n704), .A3(new_n615), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  OAI211_X1 g530(.A(new_n709), .B(new_n636), .C1(new_n599), .C2(new_n600), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n682), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n704), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  AOI21_X1  g534(.A(new_n594), .B1(new_n645), .B2(new_n537), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n379), .A2(new_n309), .A3(new_n387), .ZN(new_n722));
  AOI211_X1 g536(.A(G902), .B(new_n301), .C1(new_n652), .C2(new_n653), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n296), .A2(new_n198), .B1(new_n274), .B2(new_n277), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n268), .A2(new_n287), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n724), .A2(new_n287), .B1(new_n725), .B2(new_n650), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n290), .B1(new_n726), .B2(new_n300), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n308), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n722), .B1(new_n728), .B2(KEYINPUT102), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n308), .C1(new_n723), .C2(new_n727), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n721), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n733));
  INV_X1    g547(.A(new_n593), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n645), .B2(new_n537), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n729), .A3(new_n683), .A4(new_n731), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n732), .A2(new_n733), .B1(new_n736), .B2(KEYINPUT42), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NAND4_X1  g552(.A1(new_n721), .A2(new_n729), .A3(new_n659), .A4(new_n731), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT103), .B(G134), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G36));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n290), .B1(new_n726), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n298), .A2(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(G469), .A2(G902), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n305), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n308), .A3(new_n662), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n613), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n446), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n446), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT43), .B1(new_n758), .B2(KEYINPUT105), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n758), .B(new_n613), .C1(KEYINPUT105), .C2(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n602), .A2(new_n635), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n722), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n768), .A2(new_n769), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n772), .A2(KEYINPUT107), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT107), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n754), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n190), .ZN(G39));
  INV_X1    g591(.A(new_n556), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n595), .A2(new_n682), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n771), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n308), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT47), .B1(new_n750), .B2(new_n308), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NOR2_X1   g600(.A1(new_n695), .A2(new_n722), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n595), .A2(new_n671), .A3(new_n448), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n446), .A3(new_n613), .ZN(new_n789));
  INV_X1    g603(.A(new_n448), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n760), .B2(new_n761), .ZN(new_n791));
  INV_X1    g605(.A(new_n710), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n704), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n789), .A2(G952), .A3(new_n793), .A4(new_n391), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT48), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n791), .A2(KEYINPUT113), .A3(new_n787), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n791), .B2(new_n787), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n796), .B1(new_n799), .B2(new_n735), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n796), .A3(new_n735), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n784), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n305), .B1(new_n654), .B2(new_n290), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n803), .B(new_n782), .C1(new_n308), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n791), .A2(new_n792), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n722), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n613), .A2(new_n446), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n788), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n788), .A2(KEYINPUT114), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n717), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n797), .B2(new_n798), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n674), .A2(new_n310), .A3(new_n696), .ZN(new_n818));
  OAI211_X1 g632(.A(KEYINPUT112), .B(KEYINPUT50), .C1(new_n806), .C2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT112), .B1(new_n806), .B2(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n815), .A2(new_n817), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  OAI221_X1 g637(.A(new_n795), .B1(new_n800), .B2(new_n802), .C1(new_n809), .C2(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(KEYINPUT115), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n823), .A2(KEYINPUT115), .B1(new_n805), .B2(new_n807), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT116), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n703), .A2(new_n713), .A3(new_n712), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n636), .A2(new_n658), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n728), .A2(KEYINPUT110), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n647), .B1(new_n648), .B2(new_n305), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(new_n831), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n670), .B(new_n830), .C1(new_n833), .C2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT110), .B1(new_n728), .B2(new_n832), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n835), .A2(new_n834), .A3(new_n831), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(KEYINPUT111), .A3(new_n670), .A4(new_n830), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n660), .A2(new_n719), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n829), .A2(new_n844), .A3(new_n691), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n690), .B2(new_n685), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n829), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n697), .A2(new_n705), .A3(new_n715), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n701), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n721), .A2(new_n729), .A3(new_n659), .A4(new_n731), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n728), .A2(KEYINPUT102), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n718), .A3(new_n731), .A4(new_n771), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n497), .A2(new_n635), .A3(new_n658), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n623), .A3(new_n624), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n722), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(new_n556), .A3(new_n308), .A4(new_n306), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n499), .B1(new_n596), .B2(new_n637), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n446), .A2(new_n497), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n755), .B2(new_n446), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n388), .A3(new_n615), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n603), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n737), .A2(new_n852), .A3(new_n861), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT109), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n739), .A2(new_n855), .A3(new_n859), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n866), .A3(new_n862), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(KEYINPUT109), .A3(new_n737), .A4(new_n852), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT53), .B1(new_n845), .B2(KEYINPUT52), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n850), .B2(new_n874), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n870), .A2(new_n873), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n848), .A2(new_n844), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n848), .A2(new_n829), .A3(new_n844), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n845), .B2(KEYINPUT52), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n872), .A2(new_n888), .A3(new_n737), .A4(new_n852), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n847), .A2(new_n889), .A3(new_n849), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n828), .A2(new_n879), .A3(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT116), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n893), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n593), .A2(new_n308), .A3(new_n309), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n757), .A2(KEYINPUT108), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n674), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n804), .B(KEYINPUT49), .Z(new_n900));
  OAI21_X1  g714(.A(KEYINPUT108), .B1(new_n757), .B2(new_n896), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n671), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n902), .ZN(G75));
  INV_X1    g717(.A(new_n280), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n447), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT117), .Z(new_n906));
  AOI21_X1  g720(.A(new_n300), .B1(new_n886), .B2(new_n891), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(G210), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n348), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n385), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n906), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n910), .B2(new_n914), .ZN(G51));
  INV_X1    g730(.A(new_n745), .ZN(new_n917));
  OAI211_X1 g731(.A(G902), .B(new_n917), .C1(new_n878), .C2(new_n890), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n746), .B(KEYINPUT118), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n887), .B1(new_n886), .B2(new_n891), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n878), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n303), .A2(new_n304), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT119), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n919), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n906), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT120), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n930));
  INV_X1    g744(.A(new_n926), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n878), .B2(new_n890), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n892), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n933), .B2(new_n921), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n930), .B(new_n906), .C1(new_n934), .C2(new_n919), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n929), .A2(new_n935), .ZN(G54));
  NAND3_X1  g750(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(new_n434), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n434), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n928), .B1(new_n938), .B2(new_n939), .ZN(G60));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT59), .Z(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n879), .B2(new_n892), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n609), .A2(new_n610), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n906), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n942), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n933), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n878), .B2(new_n890), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(new_n633), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n587), .ZN(new_n955));
  NOR2_X1   g769(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n928), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT123), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n958), .B(new_n961), .ZN(G66));
  OAI21_X1  g776(.A(G953), .B1(new_n450), .B2(new_n345), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n852), .A2(new_n867), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n904), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n911), .B1(G898), .B2(new_n280), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  AOI21_X1  g781(.A(new_n280), .B1(G227), .B2(G900), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n848), .A2(new_n679), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n721), .A2(new_n771), .A3(new_n864), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n663), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT125), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n785), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n776), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n971), .A2(new_n972), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n904), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n522), .A2(new_n526), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n429), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n785), .A2(new_n737), .A3(new_n739), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n735), .A2(new_n830), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n986), .B(new_n848), .C1(new_n754), .C2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n280), .B1(new_n988), .B2(new_n776), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n904), .A2(new_n657), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT126), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n983), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n969), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(new_n991), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n984), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n968), .C1(new_n981), .C2(new_n984), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(G72));
  NAND3_X1  g811(.A1(new_n978), .A2(new_n964), .A3(new_n980), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n665), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n527), .A2(new_n529), .A3(new_n510), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n988), .A2(new_n776), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n964), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n886), .B1(new_n875), .B2(new_n876), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n530), .B1(new_n540), .B2(new_n541), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1007), .A2(new_n1000), .A3(new_n1008), .ZN(new_n1009));
  NOR4_X1   g823(.A1(new_n1002), .A2(new_n1006), .A3(new_n1009), .A4(new_n928), .ZN(G57));
endmodule


