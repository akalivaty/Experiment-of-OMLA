//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT66), .Z(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n213), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n227), .B1(new_n231), .B2(new_n233), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n223), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n215), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n259), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT69), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n228), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n271), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(G274), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n270), .B2(new_n271), .ZN(new_n281));
  XOR2_X1   g0081(.A(KEYINPUT68), .B(G226), .Z(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(G169), .ZN(new_n287));
  INV_X1    g0087(.A(G1), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT72), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n228), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n288), .A2(G13), .A3(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(new_n288), .A3(G13), .A4(G20), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n295), .A2(new_n297), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n291), .A2(new_n298), .B1(new_n202), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n293), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT8), .B(G58), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n229), .A2(G33), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n286), .A2(new_n287), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G200), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n274), .B2(new_n283), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G190), .B2(new_n284), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT9), .ZN(new_n317));
  INV_X1    g0117(.A(new_n311), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n300), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n301), .A2(new_n311), .A3(KEYINPUT9), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n316), .B(new_n323), .C1(new_n319), .C2(new_n320), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n313), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n327));
  INV_X1    g0127(.A(G107), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n327), .B1(new_n328), .B2(new_n257), .C1(new_n264), .C2(new_n216), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n329), .A2(new_n273), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n288), .B1(G41), .B2(G45), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n275), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n279), .B1(new_n332), .B2(new_n218), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n326), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G20), .A2(G77), .ZN(new_n335));
  INV_X1    g0135(.A(new_n309), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n335), .B1(new_n303), .B2(new_n336), .C1(new_n305), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n293), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n298), .A2(G77), .A3(new_n289), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n299), .A2(new_n217), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT74), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n333), .B1(new_n329), .B2(new_n273), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(KEYINPUT74), .C1(new_n344), .C2(G169), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n285), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT73), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n350), .C1(new_n314), .C2(new_n344), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n314), .B2(new_n344), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(KEYINPUT73), .B1(G190), .B2(new_n344), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  OAI211_X1 g0155(.A(G232), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n257), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n273), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n279), .B1(new_n332), .B2(new_n216), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n355), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g0166(.A(KEYINPUT13), .B(new_n364), .C1(new_n362), .C2(new_n273), .ZN(new_n367));
  OAI21_X1  g0167(.A(G200), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n299), .A2(new_n215), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT12), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n336), .A2(new_n202), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n305), .A2(new_n217), .B1(new_n229), .B2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n293), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT11), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n298), .A2(G68), .A3(new_n289), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n363), .A2(new_n365), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n363), .A2(new_n355), .A3(new_n365), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n368), .B(new_n376), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n366), .A2(new_n367), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(G190), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(KEYINPUT76), .A3(new_n368), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n380), .B2(G169), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(G169), .C1(new_n366), .C2(new_n367), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n378), .A2(G179), .A3(new_n379), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n385), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n325), .A2(new_n354), .A3(new_n389), .A4(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT7), .B1(new_n262), .B2(new_n229), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n256), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT77), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n255), .A2(new_n229), .A3(new_n256), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n215), .B1(new_n404), .B2(new_n398), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G58), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n215), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n409), .B2(new_n201), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n309), .A2(G159), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n410), .A2(KEYINPUT16), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n401), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n293), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n304), .A2(new_n307), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n288), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n298), .B1(new_n299), .B2(new_n418), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n265), .A2(new_n258), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G226), .B2(new_n258), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n422), .A2(new_n262), .B1(new_n254), .B2(new_n209), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n273), .ZN(new_n424));
  INV_X1    g0224(.A(G274), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n270), .B2(new_n271), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n281), .A2(G232), .B1(new_n278), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n427), .A3(new_n381), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n424), .A2(new_n427), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(G200), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n417), .A2(new_n420), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT17), .ZN(new_n432));
  XOR2_X1   g0232(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n417), .A2(new_n420), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n326), .B1(new_n424), .B2(new_n427), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(G179), .B2(new_n429), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n417), .B2(new_n420), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND4_X1   g0243(.A1(KEYINPUT80), .A2(new_n434), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n441), .B(KEYINPUT18), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT80), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n396), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n288), .A2(G33), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n298), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G97), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n295), .A2(new_n211), .A3(new_n297), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT82), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n328), .A2(KEYINPUT6), .A3(G97), .ZN(new_n456));
  XNOR2_X1  g0256(.A(G97), .B(G107), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT6), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n459), .A2(new_n229), .B1(new_n217), .B2(new_n336), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n328), .B1(new_n404), .B2(new_n398), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n293), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n463));
  OAI21_X1  g0263(.A(G107), .B1(new_n397), .B2(new_n399), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n336), .A2(new_n217), .ZN(new_n465));
  AND2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n328), .A2(KEYINPUT6), .A3(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n470), .B2(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT81), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(new_n293), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n455), .B1(new_n463), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n273), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n288), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT83), .A3(new_n288), .A4(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n487), .A2(G41), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n486), .A2(new_n489), .A3(new_n426), .A4(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n275), .B(G257), .C1(new_n484), .C2(new_n490), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(KEYINPUT84), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n483), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G190), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n492), .A2(KEYINPUT84), .A3(new_n493), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT84), .B1(new_n492), .B2(new_n493), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(G200), .B1(new_n502), .B2(new_n483), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n475), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n451), .A2(new_n454), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n473), .B1(new_n472), .B2(new_n293), .ZN(new_n506));
  AOI211_X1 g0306(.A(KEYINPUT81), .B(new_n302), .C1(new_n464), .C2(new_n471), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n285), .A3(new_n483), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n498), .A2(new_n326), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n229), .B1(new_n512), .B2(new_n360), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n467), .A2(new_n209), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(new_n255), .B2(new_n256), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n229), .A2(G33), .A3(G97), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n516), .A2(G68), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n293), .B1(new_n299), .B2(new_n337), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n298), .A2(G87), .A3(new_n449), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT86), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n298), .A2(KEYINPUT86), .A3(G87), .A4(new_n449), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n288), .A2(new_n425), .A3(G45), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n210), .B1(new_n277), .B2(G1), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n275), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n530));
  OAI211_X1 g0330(.A(G238), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n531));
  INV_X1    g0331(.A(G116), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n254), .C2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n381), .B(new_n529), .C1(new_n533), .C2(new_n273), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n529), .B1(new_n533), .B2(new_n273), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n534), .B1(G200), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n535), .A2(G169), .ZN(new_n538));
  AOI211_X1 g0338(.A(G179), .B(new_n529), .C1(new_n533), .C2(new_n273), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n519), .A2(new_n293), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n299), .A2(new_n337), .ZN(new_n542));
  INV_X1    g0342(.A(new_n337), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n450), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n526), .A2(new_n537), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n504), .A2(new_n511), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n298), .A2(G116), .A3(new_n449), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n299), .A2(new_n532), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n292), .A2(new_n228), .B1(G20), .B2(new_n532), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n480), .B(new_n229), .C1(G33), .C2(new_n211), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n552), .A2(KEYINPUT20), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT20), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n255), .A2(G303), .A3(new_n256), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n273), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n275), .B(G270), .C1(new_n484), .C2(new_n490), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(G179), .A3(new_n492), .A4(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n548), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  AND4_X1   g0365(.A1(G179), .A2(new_n562), .A3(new_n492), .A4(new_n563), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n549), .B(new_n550), .C1(new_n555), .C2(new_n554), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(KEYINPUT87), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n492), .A3(new_n563), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(G169), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n567), .A2(KEYINPUT21), .A3(new_n570), .A4(G169), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(G200), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(new_n557), .C1(new_n381), .C2(new_n570), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n569), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n229), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n578));
  NAND2_X1  g0378(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n257), .A2(new_n229), .A3(G87), .A4(new_n579), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n229), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n328), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n306), .A2(G116), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n584), .B1(new_n583), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n293), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n328), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n295), .A2(new_n297), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(G107), .ZN(new_n595));
  AOI22_X1  g0395(.A1(G107), .A2(new_n450), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n275), .B(G264), .C1(new_n484), .C2(new_n490), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G250), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n212), .B2(G1698), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n257), .B1(G33), .B2(G294), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n269), .A2(new_n272), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(KEYINPUT89), .B(new_n598), .C1(new_n601), .C2(new_n602), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(G179), .A3(new_n492), .A4(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n492), .B(new_n598), .C1(new_n601), .C2(new_n602), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G169), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n597), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n608), .A2(G190), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n492), .A3(new_n606), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n314), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n597), .B2(new_n614), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n448), .A2(new_n547), .A3(new_n577), .A4(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n347), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT74), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n344), .A2(G169), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n349), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n384), .B2(new_n388), .ZN(new_n622));
  INV_X1    g0422(.A(new_n395), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n434), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n445), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n322), .A2(new_n324), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n313), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n573), .A2(new_n574), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n597), .A2(new_n610), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n597), .B2(new_n610), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n569), .B(new_n628), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n504), .A2(new_n511), .A3(new_n546), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n614), .A2(new_n597), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n538), .ZN(new_n637));
  INV_X1    g0437(.A(new_n539), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n545), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n536), .A2(G200), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n535), .A2(G190), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n642), .A2(new_n520), .A3(new_n525), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n641), .B1(new_n511), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(G169), .B1(new_n502), .B2(new_n483), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n285), .A2(new_n483), .A3(new_n496), .A4(new_n497), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n546), .A2(KEYINPUT26), .A3(new_n508), .A4(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n640), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n627), .B1(new_n448), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT91), .Z(G369));
  NAND3_X1  g0455(.A1(new_n288), .A2(new_n229), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT92), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(G343), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(G343), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n567), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n628), .A2(new_n569), .A3(new_n576), .A4(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n628), .A2(new_n569), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT93), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT93), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n670), .A3(G330), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n597), .A2(new_n663), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT94), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n597), .A2(KEYINPUT94), .A3(new_n663), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n635), .A2(new_n675), .A3(new_n611), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n597), .A2(new_n610), .A3(new_n663), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT95), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT95), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n597), .A2(new_n610), .A3(new_n680), .A4(new_n663), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT96), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n677), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n672), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n630), .A2(new_n631), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n663), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n666), .A2(new_n663), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n224), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n514), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n233), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n504), .A2(new_n511), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n628), .A2(new_n569), .A3(new_n611), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n546), .A3(new_n703), .A4(new_n635), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n651), .ZN(new_n705));
  INV_X1    g0505(.A(new_n663), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI211_X1 g0507(.A(KEYINPUT29), .B(new_n663), .C1(new_n636), .C2(new_n651), .ZN(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n566), .A2(new_n535), .A3(new_n605), .A4(new_n606), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n498), .ZN(new_n712));
  INV_X1    g0512(.A(new_n498), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n605), .A2(new_n535), .A3(new_n606), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(KEYINPUT30), .A4(new_n566), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n570), .A2(new_n285), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n613), .A3(new_n498), .A4(new_n536), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT31), .B1(new_n718), .B2(new_n663), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n615), .A2(new_n577), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n633), .A3(new_n706), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n709), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NOR4_X1   g0524(.A1(new_n707), .A2(new_n708), .A3(new_n724), .A4(KEYINPUT97), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT97), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n708), .A2(new_n707), .ZN(new_n727));
  INV_X1    g0527(.A(new_n724), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n700), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n672), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n229), .A2(G13), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n288), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n695), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n733), .B(new_n739), .C1(G330), .C2(new_n667), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n228), .B1(G20), .B2(new_n326), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT99), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n251), .A2(new_n277), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n694), .A2(new_n257), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G45), .B2(new_n233), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n257), .A2(new_n224), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n224), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n751), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n746), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n229), .A2(new_n285), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n381), .A3(G200), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT33), .B(G317), .Z(new_n760));
  NOR2_X1   g0560(.A1(new_n229), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n381), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n759), .A2(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n257), .B1(new_n767), .B2(G329), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n758), .A2(new_n765), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n381), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n764), .B(new_n771), .C1(G322), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n758), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n381), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n780), .A2(G326), .B1(new_n782), .B2(G303), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n285), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n778), .B(new_n783), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n789));
  INV_X1    g0589(.A(new_n780), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n767), .A2(G159), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n790), .A2(new_n202), .B1(new_n791), .B2(KEYINPUT32), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n759), .A2(new_n215), .B1(new_n762), .B2(new_n328), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n777), .A2(G58), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n257), .B1(new_n770), .B2(new_n217), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(KEYINPUT32), .B2(new_n791), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n782), .A2(G87), .B1(new_n786), .B2(G97), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n794), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n789), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n739), .B(new_n757), .C1(new_n801), .C2(new_n744), .ZN(new_n802));
  INV_X1    g0602(.A(new_n743), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n667), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n740), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n349), .A2(new_n706), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n353), .B2(new_n351), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT104), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n343), .B2(new_n347), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n617), .A2(KEYINPUT104), .A3(new_n620), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n348), .A2(new_n807), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n724), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n718), .A2(new_n663), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT31), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n547), .A2(new_n615), .A3(new_n577), .A4(new_n663), .ZN(new_n821));
  OAI211_X1 g0621(.A(G330), .B(new_n814), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n663), .B1(new_n636), .B2(new_n651), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n815), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n815), .B2(new_n823), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n738), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n814), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n741), .ZN(new_n831));
  INV_X1    g0631(.A(new_n759), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(G150), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n770), .C1(new_n790), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G143), .B2(new_n777), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n257), .B1(new_n766), .B2(new_n839), .C1(new_n787), .C2(new_n408), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n202), .A2(new_n781), .B1(new_n762), .B2(new_n215), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G303), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n790), .A2(new_n843), .B1(new_n770), .B2(new_n532), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G283), .B2(new_n832), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT102), .Z(new_n846));
  AOI22_X1  g0646(.A1(new_n777), .A2(G294), .B1(G97), .B2(new_n786), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n262), .B1(new_n766), .B2(new_n769), .C1(new_n328), .C2(new_n781), .ZN(new_n850));
  INV_X1    g0650(.A(new_n762), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(G87), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n838), .A2(new_n842), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n744), .A2(new_n741), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n854), .A2(new_n744), .B1(new_n217), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n739), .B1(new_n831), .B2(new_n856), .ZN(new_n857));
  OR3_X1    g0657(.A1(new_n829), .A2(KEYINPUT105), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT105), .B1(new_n829), .B2(new_n857), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  AOI211_X1 g0661(.A(new_n532), .B(new_n231), .C1(new_n470), .C2(KEYINPUT35), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(KEYINPUT35), .B2(new_n470), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT36), .Z(new_n864));
  OR3_X1    g0664(.A1(new_n233), .A2(new_n217), .A3(new_n409), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n288), .B(G13), .C1(new_n865), .C2(new_n247), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n419), .A2(new_n298), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n418), .A2(new_n299), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n413), .A2(new_n293), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n401), .A2(new_n407), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n414), .B1(new_n873), .B2(new_n415), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n431), .B1(new_n875), .B2(new_n659), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n437), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n659), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n435), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n439), .A2(new_n880), .A3(new_n881), .A4(new_n431), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(KEYINPUT107), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n434), .A2(new_n440), .A3(new_n443), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n875), .A2(new_n659), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT107), .B1(new_n878), .B2(new_n882), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n878), .A2(new_n882), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT107), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n892), .A2(KEYINPUT38), .A3(new_n886), .A4(new_n883), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n721), .A2(new_n723), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n814), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n385), .A2(new_n663), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n389), .A2(new_n395), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n389), .B2(new_n395), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n887), .A2(new_n888), .ZN(new_n905));
  INV_X1    g0705(.A(new_n880), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n439), .A2(new_n880), .A3(new_n431), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n884), .A2(new_n906), .B1(new_n908), .B2(new_n882), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT108), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT108), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n882), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n880), .B1(new_n445), .B2(new_n434), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n911), .B(new_n868), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n905), .A2(KEYINPUT38), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n382), .A2(new_n383), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT76), .B1(new_n387), .B2(new_n368), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n395), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n897), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n389), .A2(new_n395), .A3(new_n897), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n923), .A2(new_n895), .A3(KEYINPUT40), .A4(new_n814), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n904), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n447), .A2(new_n895), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(G330), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n623), .A2(new_n706), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(new_n916), .C2(KEYINPUT39), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n445), .A2(new_n879), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n824), .A2(new_n814), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n811), .A2(new_n810), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n706), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(KEYINPUT106), .A3(new_n706), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n900), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n934), .B1(new_n894), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n447), .B1(new_n708), .B2(new_n707), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n627), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n929), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n288), .B2(new_n735), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n929), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n867), .B1(new_n949), .B2(new_n950), .ZN(G367));
  OAI21_X1  g0751(.A(new_n702), .B1(new_n475), .B2(new_n706), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n649), .A2(new_n508), .A3(new_n663), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n688), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT111), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n952), .A2(new_n611), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n663), .B1(new_n958), .B2(new_n511), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n687), .A2(new_n691), .A3(new_n954), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(KEYINPUT42), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n677), .A2(new_n685), .A3(new_n682), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n685), .B1(new_n677), .B2(new_n682), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n691), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n964), .A2(KEYINPUT42), .A3(new_n955), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n526), .A2(new_n706), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n640), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n645), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(KEYINPUT110), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT109), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(KEYINPUT110), .B2(new_n970), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n966), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n972), .B1(new_n966), .B2(new_n975), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n957), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n966), .A2(new_n975), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n971), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT111), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n956), .B(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n966), .A2(new_n972), .A3(new_n975), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n695), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n692), .B2(new_n954), .ZN(new_n988));
  INV_X1    g0788(.A(new_n690), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n964), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n990), .B2(new_n955), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n954), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n688), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n992), .A2(new_n996), .A3(new_n688), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n684), .B(new_n686), .C1(new_n666), .C2(new_n663), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n964), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT112), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n733), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n964), .B(new_n1001), .C1(new_n672), .C2(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n729), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n725), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n999), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n986), .B1(new_n1010), .B2(new_n731), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n985), .B1(new_n1011), .B2(new_n737), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n748), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n745), .B1(new_n224), .B2(new_n337), .C1(new_n242), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n738), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n781), .A2(new_n532), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT46), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n777), .B2(G303), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G294), .A2(new_n832), .B1(new_n851), .B2(G97), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n780), .A2(G311), .B1(new_n786), .B2(G107), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n262), .B1(new_n766), .B2(new_n1021), .C1(new_n763), .C2(new_n770), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT46), .B2(new_n1016), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n257), .B1(new_n770), .B2(new_n202), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G137), .B2(new_n767), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G159), .A2(new_n832), .B1(new_n851), .B2(G77), .ZN(new_n1027));
  INV_X1    g0827(.A(G150), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1027), .C1(new_n1028), .C2(new_n776), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n787), .A2(new_n215), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G143), .B2(new_n780), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n408), .B2(new_n781), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1015), .B1(new_n1034), .B2(new_n744), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n969), .A2(new_n803), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1012), .A2(new_n1037), .ZN(G387));
  OAI22_X1  g0838(.A1(new_n752), .A2(new_n697), .B1(G107), .B2(new_n224), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n239), .A2(new_n277), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n697), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G45), .B(new_n1041), .C1(G68), .C2(G77), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n303), .A2(G50), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1013), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n746), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n739), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n257), .B1(new_n770), .B2(new_n215), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G150), .B2(new_n767), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n418), .B2(new_n759), .C1(new_n202), .C2(new_n776), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n217), .A2(new_n781), .B1(new_n762), .B2(new_n211), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n787), .A2(new_n337), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n790), .A2(new_n834), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n759), .A2(new_n769), .B1(new_n770), .B2(new_n843), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G322), .B2(new_n780), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1021), .B2(new_n776), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n782), .A2(G294), .B1(new_n786), .B2(G283), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT49), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT114), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n257), .B1(new_n767), .B2(G326), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n532), .B2(new_n762), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1056), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT115), .Z(new_n1073));
  INV_X1    g0873(.A(new_n744), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1049), .B1(new_n687), .B2(new_n803), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1004), .A2(new_n737), .A3(new_n1005), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n730), .A2(new_n1006), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1005), .B(new_n1004), .C1(new_n725), .C2(new_n729), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n695), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(G393));
  AND3_X1   g0881(.A1(new_n992), .A2(new_n996), .A3(new_n688), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n688), .B1(new_n992), .B2(new_n996), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n1010), .A3(new_n695), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n955), .A2(new_n743), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n745), .B1(new_n211), .B2(new_n224), .C1(new_n246), .C2(new_n1013), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n738), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n776), .A2(new_n834), .B1(new_n1028), .B2(new_n790), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT51), .Z(new_n1091));
  NOR2_X1   g0891(.A1(new_n787), .A2(new_n217), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G68), .B2(new_n782), .ZN(new_n1093));
  INV_X1    g0893(.A(G143), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n257), .B1(new_n766), .B2(new_n1094), .C1(new_n303), .C2(new_n770), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G50), .A2(new_n832), .B1(new_n851), .B2(G87), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n776), .A2(new_n769), .B1(new_n1021), .B2(new_n790), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  OAI21_X1  g0900(.A(new_n262), .B1(new_n770), .B2(new_n784), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G322), .B2(new_n767), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G303), .A2(new_n832), .B1(new_n851), .B2(G107), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n782), .A2(G283), .B1(new_n786), .B2(G116), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1091), .A2(new_n1098), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1089), .B1(new_n1106), .B2(new_n744), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1086), .A2(new_n737), .B1(new_n1087), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1085), .A2(new_n1108), .ZN(G390));
  NAND2_X1  g0909(.A1(new_n884), .A2(new_n906), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n912), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n911), .B1(new_n1111), .B2(new_n868), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n909), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n893), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT39), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n742), .B1(new_n1116), .B2(new_n932), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n739), .B1(new_n418), .B2(new_n855), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT53), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n782), .A2(new_n1119), .A3(G150), .ZN(new_n1120));
  OAI21_X1  g0920(.A(KEYINPUT53), .B1(new_n781), .B2(new_n1028), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n262), .B1(new_n767), .B2(G125), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n770), .B2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1122), .B(new_n1125), .C1(G132), .C2(new_n777), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n759), .A2(new_n835), .B1(new_n762), .B2(new_n202), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n787), .A2(new_n834), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(G128), .C2(new_n780), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n759), .A2(new_n328), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1130), .B(new_n1092), .C1(G283), .C2(new_n780), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n262), .B1(new_n766), .B2(new_n784), .C1(new_n211), .C2(new_n770), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n215), .A2(new_n762), .B1(new_n781), .B2(new_n209), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(new_n777), .C2(G116), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1126), .A2(new_n1129), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1118), .B1(new_n1135), .B2(new_n1074), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1117), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n939), .A2(new_n940), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n824), .B2(new_n814), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n930), .B1(new_n1139), .B2(new_n900), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n910), .A2(new_n915), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT39), .B1(new_n1141), .B2(new_n893), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n889), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n724), .A2(new_n814), .A3(new_n923), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n663), .B1(new_n704), .B2(new_n651), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n814), .B1(new_n706), .B2(new_n936), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1114), .B(new_n930), .C1(new_n900), .C2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1137), .B1(new_n1151), .B2(new_n737), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n935), .A2(new_n941), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n923), .B1(new_n724), .B2(new_n814), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n822), .A2(new_n900), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n822), .A2(new_n900), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1145), .A2(new_n1157), .A3(new_n1147), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n447), .A2(new_n724), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n945), .A2(new_n627), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT116), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT116), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n945), .A2(new_n1163), .A3(new_n627), .A4(new_n1160), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1159), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n695), .B1(new_n1151), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n942), .A2(new_n931), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1116), .B2(new_n932), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1147), .A2(new_n900), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n916), .A2(new_n931), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1155), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1144), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n1165), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1152), .B1(new_n1166), .B2(new_n1174), .ZN(G378));
  AOI211_X1 g0975(.A(G41), .B(new_n257), .C1(new_n767), .C2(G283), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n337), .B2(new_n770), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1030), .B(new_n1177), .C1(G77), .C2(new_n782), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n759), .A2(new_n211), .B1(new_n762), .B2(new_n408), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G116), .B2(new_n780), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n328), .C2(new_n776), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT58), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT58), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n254), .A2(new_n276), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT117), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G50), .B(new_n1186), .C1(new_n276), .C2(new_n262), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n759), .A2(new_n839), .B1(new_n770), .B2(new_n835), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n777), .B2(G128), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n780), .A2(G125), .B1(new_n786), .B2(G150), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n781), .C2(new_n1124), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n767), .A2(G124), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n1186), .C1(new_n834), .C2(new_n762), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1191), .B2(KEYINPUT59), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1187), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1183), .A2(new_n1184), .A3(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(new_n744), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n739), .B(new_n1198), .C1(new_n202), .C2(new_n855), .ZN(new_n1199));
  XOR2_X1   g0999(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n312), .A2(new_n659), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n322), .A2(new_n324), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n313), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT119), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n325), .B1(new_n312), .B2(new_n659), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1205), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1201), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1209), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n741), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1199), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(G330), .B1(new_n916), .B2(new_n924), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT40), .B1(new_n894), .B2(new_n901), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n924), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n709), .B1(new_n1114), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n904), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n944), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n904), .A2(new_n1221), .A3(new_n1213), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n933), .A4(new_n943), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1215), .B1(new_n1227), .B2(new_n736), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1151), .B2(new_n1159), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1223), .A2(new_n1226), .A3(KEYINPUT57), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n695), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1230), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1173), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1229), .B1(new_n1233), .B2(new_n1237), .ZN(G375));
  AND2_X1   g1038(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1230), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n986), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1159), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n790), .A2(new_n839), .B1(new_n781), .B2(new_n834), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G50), .B2(new_n786), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n777), .A2(G137), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n770), .A2(new_n1028), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n262), .B(new_n1247), .C1(G128), .C2(new_n767), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1124), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n832), .A2(new_n1249), .B1(new_n851), .B2(G58), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n777), .A2(G283), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1054), .B1(G77), .B2(new_n851), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n759), .A2(new_n532), .B1(new_n781), .B2(new_n211), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G294), .B2(new_n780), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n262), .B1(new_n770), .B2(new_n328), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G303), .B2(new_n767), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1252), .A2(new_n1253), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1074), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n739), .B(new_n1259), .C1(new_n215), .C2(new_n855), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n923), .B2(new_n742), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1239), .B2(new_n736), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1243), .A2(new_n1263), .ZN(G381));
  NAND3_X1  g1064(.A1(new_n1077), .A2(new_n1080), .A3(new_n805), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G384), .A2(G390), .A3(new_n1265), .A4(G381), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(new_n1266), .A2(G375), .A3(G387), .A4(G378), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT120), .Z(G407));
  NAND2_X1  g1068(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1269), .A2(new_n736), .B1(new_n1117), .B2(new_n1136), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n696), .B1(new_n1269), .B2(new_n1242), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1173), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n661), .A2(new_n662), .A3(G213), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G375), .C2(new_n1275), .ZN(G409));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  INV_X1    g1077(.A(G390), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n978), .A2(new_n984), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1082), .A2(new_n1083), .A3(new_n1079), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1241), .B1(new_n1280), .B2(new_n730), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1281), .B2(new_n736), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1037), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1012), .A2(new_n1037), .A3(G390), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1265), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G390), .B1(new_n1012), .B2(new_n1037), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(KEYINPUT124), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(new_n1286), .A3(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT125), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1284), .A2(new_n1295), .A3(new_n1286), .A4(new_n1289), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1274), .A2(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT121), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1159), .B1(new_n1164), .B2(new_n1162), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n695), .B1(new_n1302), .B2(KEYINPUT60), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1299), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT60), .B1(new_n1165), .B2(new_n1302), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n696), .B1(new_n1240), .B2(new_n1300), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(KEYINPUT121), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G384), .B1(new_n1308), .B2(new_n1263), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n860), .B(new_n1262), .C1(new_n1304), .C2(new_n1307), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1274), .A2(KEYINPUT123), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1298), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1301), .A2(new_n1303), .A3(new_n1299), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT121), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1263), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n860), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1308), .A2(G384), .A3(new_n1263), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1317), .A2(new_n1298), .A3(new_n1318), .A4(new_n1312), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1313), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G378), .B(new_n1229), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1234), .A2(new_n1236), .A3(new_n1241), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1272), .B1(new_n1323), .B2(new_n1228), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1273), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1321), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1274), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1311), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1328), .B2(new_n1311), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1297), .B1(new_n1327), .B2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1325), .A2(new_n1273), .A3(new_n1311), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1311), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1336), .A2(new_n1297), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1317), .A2(new_n1318), .A3(new_n1312), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1298), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1319), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT122), .B1(new_n1325), .B2(new_n1273), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT122), .ZN(new_n1345));
  AOI211_X1 g1145(.A(new_n1345), .B(new_n1274), .C1(new_n1322), .C2(new_n1324), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1343), .A2(new_n1344), .A3(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1339), .A2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1277), .B1(new_n1333), .B2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1326), .A2(new_n1342), .A3(new_n1319), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1334), .A2(KEYINPUT62), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1328), .A2(new_n1329), .A3(new_n1311), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1350), .A2(new_n1351), .A3(new_n1337), .A4(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1297), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1355), .B(KEYINPUT126), .C1(new_n1347), .C2(new_n1339), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1349), .A2(new_n1356), .ZN(G405));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1272), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1359), .A2(new_n1322), .A3(new_n1311), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1311), .B1(new_n1359), .B2(new_n1322), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1358), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1297), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1360), .A2(new_n1361), .A3(new_n1358), .ZN(new_n1364));
  XNOR2_X1  g1164(.A(new_n1363), .B(new_n1364), .ZN(G402));
endmodule


