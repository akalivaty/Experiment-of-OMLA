

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U550 ( .A1(n726), .A2(n725), .ZN(n777) );
  AND2_X1 U551 ( .A1(n554), .A2(G2104), .ZN(n894) );
  NOR2_X4 U552 ( .A1(n798), .A2(n688), .ZN(n725) );
  XNOR2_X2 U553 ( .A(KEYINPUT71), .B(n587), .ZN(n1019) );
  BUF_X1 U554 ( .A(n685), .Z(G160) );
  BUF_X1 U555 ( .A(n620), .Z(n621) );
  XNOR2_X1 U556 ( .A(n722), .B(n721), .ZN(n723) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n721) );
  XNOR2_X1 U558 ( .A(n582), .B(KEYINPUT13), .ZN(n583) );
  XNOR2_X1 U559 ( .A(n774), .B(KEYINPUT99), .ZN(n778) );
  XOR2_X1 U560 ( .A(KEYINPUT66), .B(G651), .Z(n519) );
  NOR2_X1 U561 ( .A1(n765), .A2(n777), .ZN(n520) );
  AND2_X1 U562 ( .A1(n553), .A2(n552), .ZN(n521) );
  NAND2_X1 U563 ( .A1(n744), .A2(G303), .ZN(n522) );
  NOR2_X1 U564 ( .A1(n766), .A2(n777), .ZN(n523) );
  AND2_X1 U565 ( .A1(n731), .A2(n730), .ZN(n524) );
  OR2_X1 U566 ( .A1(n777), .A2(n776), .ZN(n525) );
  AND2_X1 U567 ( .A1(n710), .A2(n709), .ZN(n526) );
  AND2_X1 U568 ( .A1(n711), .A2(n526), .ZN(n712) );
  NOR2_X1 U569 ( .A1(n713), .A2(n712), .ZN(n714) );
  INV_X1 U570 ( .A(KEYINPUT31), .ZN(n734) );
  XNOR2_X1 U571 ( .A(n734), .B(KEYINPUT96), .ZN(n735) );
  XNOR2_X1 U572 ( .A(n736), .B(n735), .ZN(n737) );
  INV_X1 U573 ( .A(KEYINPUT97), .ZN(n739) );
  INV_X1 U574 ( .A(KEYINPUT70), .ZN(n582) );
  NOR2_X1 U575 ( .A1(G164), .A2(G1384), .ZN(n687) );
  AND2_X1 U576 ( .A1(n778), .A2(n525), .ZN(n779) );
  XNOR2_X1 U577 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n551) );
  NOR2_X1 U579 ( .A1(n639), .A2(n519), .ZN(n647) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U581 ( .A1(n649), .A2(G89), .ZN(n527) );
  XNOR2_X1 U582 ( .A(n527), .B(KEYINPUT4), .ZN(n529) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  NAND2_X1 U584 ( .A1(G76), .A2(n647), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n530), .B(KEYINPUT5), .ZN(n536) );
  NOR2_X1 U587 ( .A1(G651), .A2(n639), .ZN(n650) );
  NAND2_X1 U588 ( .A1(n650), .A2(G51), .ZN(n533) );
  NOR2_X1 U589 ( .A1(G543), .A2(n519), .ZN(n531) );
  XOR2_X2 U590 ( .A(KEYINPUT1), .B(n531), .Z(n653) );
  NAND2_X1 U591 ( .A1(G63), .A2(n653), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U593 ( .A(KEYINPUT6), .B(n534), .Z(n535) );
  NAND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U596 ( .A1(G90), .A2(n649), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G77), .A2(n647), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U599 ( .A(KEYINPUT9), .B(n540), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n653), .A2(G64), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n650), .A2(G52), .ZN(n541) );
  AND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(G301) );
  INV_X1 U604 ( .A(G301), .ZN(G171) );
  NAND2_X1 U605 ( .A1(n650), .A2(G47), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G60), .A2(n653), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G85), .A2(n649), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G72), .A2(n647), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U611 ( .A1(n550), .A2(n549), .ZN(G290) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U613 ( .A(KEYINPUT17), .B(n551), .Z(n620) );
  AND2_X1 U614 ( .A1(n620), .A2(G138), .ZN(n557) );
  INV_X1 U615 ( .A(G2105), .ZN(n554) );
  NOR2_X1 U616 ( .A1(G2104), .A2(n554), .ZN(n616) );
  NAND2_X1 U617 ( .A1(G126), .A2(n616), .ZN(n553) );
  AND2_X1 U618 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U619 ( .A1(G114), .A2(n898), .ZN(n552) );
  NAND2_X1 U620 ( .A1(G102), .A2(n894), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n521), .A2(n555), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(G164) );
  BUF_X1 U623 ( .A(n616), .Z(n873) );
  NAND2_X1 U624 ( .A1(G125), .A2(n873), .ZN(n559) );
  NAND2_X1 U625 ( .A1(G137), .A2(n620), .ZN(n558) );
  AND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G101), .A2(n894), .ZN(n560) );
  XNOR2_X1 U628 ( .A(KEYINPUT23), .B(n560), .ZN(n562) );
  AND2_X1 U629 ( .A1(n898), .A2(G113), .ZN(n561) );
  NOR2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT65), .ZN(n685) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G82), .ZN(G220) );
  NAND2_X1 U636 ( .A1(n650), .A2(G50), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G62), .A2(n653), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G88), .A2(n649), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G75), .A2(n647), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT78), .B(n573), .Z(G303) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U645 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U646 ( .A(G223), .ZN(n833) );
  NAND2_X1 U647 ( .A1(n833), .A2(G567), .ZN(n575) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U649 ( .A1(G56), .A2(n653), .ZN(n576) );
  XNOR2_X1 U650 ( .A(n576), .B(KEYINPUT14), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G43), .A2(n650), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n649), .A2(G81), .ZN(n579) );
  XNOR2_X1 U654 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G68), .A2(n647), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U658 ( .A(n1019), .ZN(n612) );
  NAND2_X1 U659 ( .A1(n612), .A2(G860), .ZN(G153) );
  NAND2_X1 U660 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G92), .A2(n649), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G79), .A2(n647), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n650), .A2(G54), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G66), .A2(n653), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U668 ( .A(n594), .B(KEYINPUT15), .ZN(n708) );
  INV_X1 U669 ( .A(n708), .ZN(n595) );
  INV_X1 U670 ( .A(n595), .ZN(n1007) );
  INV_X1 U671 ( .A(G868), .ZN(n668) );
  NAND2_X1 U672 ( .A1(n1007), .A2(n668), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(G284) );
  XOR2_X1 U674 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U675 ( .A1(n647), .A2(G78), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT67), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n650), .A2(G53), .ZN(n599) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT68), .ZN(n601) );
  NAND2_X1 U679 ( .A1(G65), .A2(n653), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U681 ( .A(KEYINPUT69), .B(n602), .Z(n603) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n649), .A2(G91), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(G299) );
  NOR2_X1 U685 ( .A1(G286), .A2(n668), .ZN(n608) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(G297) );
  INV_X1 U688 ( .A(G860), .ZN(n630) );
  NAND2_X1 U689 ( .A1(n630), .A2(G559), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n609), .A2(n595), .ZN(n610) );
  XNOR2_X1 U691 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G559), .A2(n1007), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n668), .A2(n611), .ZN(n614) );
  NOR2_X1 U694 ( .A1(n612), .A2(G868), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U696 ( .A(KEYINPUT72), .B(n615), .Z(G282) );
  NAND2_X1 U697 ( .A1(n616), .A2(G123), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n617), .B(KEYINPUT18), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G111), .A2(n898), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G99), .A2(n894), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G135), .A2(n621), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n974) );
  XNOR2_X1 U705 ( .A(G2096), .B(n974), .ZN(n627) );
  INV_X1 U706 ( .A(G2100), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(G156) );
  XNOR2_X1 U708 ( .A(n1019), .B(KEYINPUT73), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n595), .A2(G559), .ZN(n628) );
  XNOR2_X1 U710 ( .A(n629), .B(n628), .ZN(n666) );
  NAND2_X1 U711 ( .A1(n630), .A2(n666), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n650), .A2(G55), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G67), .A2(n653), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n649), .A2(G93), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT74), .B(n633), .Z(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G80), .A2(n647), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n669) );
  XNOR2_X1 U720 ( .A(n638), .B(n669), .ZN(G145) );
  NAND2_X1 U721 ( .A1(G87), .A2(n639), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G49), .A2(n650), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U725 ( .A1(n653), .A2(n642), .ZN(n643) );
  XOR2_X1 U726 ( .A(KEYINPUT75), .B(n643), .Z(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U728 ( .A(n646), .B(KEYINPUT76), .ZN(G288) );
  NAND2_X1 U729 ( .A1(n647), .A2(G73), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(KEYINPUT2), .ZN(n658) );
  NAND2_X1 U731 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G48), .A2(n650), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U734 ( .A1(G61), .A2(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(KEYINPUT77), .B(n654), .ZN(n655) );
  NOR2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(G305) );
  INV_X1 U738 ( .A(G299), .ZN(n716) );
  XNOR2_X1 U739 ( .A(n716), .B(G288), .ZN(n665) );
  XNOR2_X1 U740 ( .A(G303), .B(n669), .ZN(n662) );
  XNOR2_X1 U741 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n660) );
  XNOR2_X1 U742 ( .A(G305), .B(KEYINPUT19), .ZN(n659) );
  XNOR2_X1 U743 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n663), .B(G290), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n665), .B(n664), .ZN(n859) );
  XNOR2_X1 U747 ( .A(n666), .B(n859), .ZN(n667) );
  NOR2_X1 U748 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U749 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U750 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n675), .A2(G2072), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT81), .B(n676), .Z(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G96), .A2(n679), .ZN(n837) );
  NAND2_X1 U762 ( .A1(n837), .A2(G2106), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U764 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U765 ( .A1(G108), .A2(n681), .ZN(n838) );
  NAND2_X1 U766 ( .A1(n838), .A2(G567), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n839) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U769 ( .A1(n839), .A2(n684), .ZN(n836) );
  NAND2_X1 U770 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U771 ( .A1(n685), .A2(G40), .ZN(n798) );
  XNOR2_X1 U772 ( .A(n687), .B(KEYINPUT64), .ZN(n797) );
  INV_X1 U773 ( .A(n797), .ZN(n688) );
  XNOR2_X1 U774 ( .A(KEYINPUT25), .B(G2078), .ZN(n951) );
  NAND2_X1 U775 ( .A1(n725), .A2(n951), .ZN(n689) );
  XOR2_X1 U776 ( .A(KEYINPUT88), .B(n689), .Z(n691) );
  NOR2_X1 U777 ( .A1(n725), .A2(G1961), .ZN(n690) );
  NOR2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U779 ( .A(KEYINPUT89), .B(n692), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G171), .ZN(n724) );
  INV_X1 U781 ( .A(n725), .ZN(n741) );
  NAND2_X1 U782 ( .A1(G1956), .A2(n741), .ZN(n695) );
  NAND2_X1 U783 ( .A1(n725), .A2(G2072), .ZN(n693) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(n693), .Z(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT90), .B(n696), .Z(n715) );
  NOR2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n698) );
  XNOR2_X1 U788 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n697) );
  XNOR2_X1 U789 ( .A(n698), .B(n697), .ZN(n720) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n741), .ZN(n700) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n725), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n707) );
  NOR2_X1 U793 ( .A1(n1007), .A2(n707), .ZN(n713) );
  INV_X1 U794 ( .A(G1341), .ZN(n701) );
  OR2_X1 U795 ( .A1(n701), .A2(n725), .ZN(n702) );
  XNOR2_X1 U796 ( .A(KEYINPUT93), .B(n702), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n1019), .A2(n703), .ZN(n711) );
  XOR2_X1 U798 ( .A(KEYINPUT26), .B(KEYINPUT92), .Z(n705) );
  NAND2_X1 U799 ( .A1(n725), .A2(G1996), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n705), .B(n704), .ZN(n706) );
  INV_X1 U801 ( .A(n706), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U803 ( .A(n714), .B(KEYINPUT94), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U807 ( .A1(n724), .A2(n723), .ZN(n738) );
  INV_X1 U808 ( .A(G8), .ZN(n726) );
  NOR2_X1 U809 ( .A1(G1966), .A2(n777), .ZN(n751) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n741), .ZN(n748) );
  NOR2_X1 U811 ( .A1(n751), .A2(n748), .ZN(n727) );
  NAND2_X1 U812 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U813 ( .A(n728), .B(KEYINPUT30), .ZN(n729) );
  XNOR2_X1 U814 ( .A(n729), .B(KEYINPUT95), .ZN(n731) );
  INV_X1 U815 ( .A(G168), .ZN(n730) );
  NOR2_X1 U816 ( .A1(G171), .A2(n732), .ZN(n733) );
  NOR2_X1 U817 ( .A1(n524), .A2(n733), .ZN(n736) );
  NAND2_X1 U818 ( .A1(n738), .A2(n737), .ZN(n749) );
  NAND2_X1 U819 ( .A1(G286), .A2(n749), .ZN(n740) );
  XNOR2_X1 U820 ( .A(n740), .B(n739), .ZN(n745) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n777), .ZN(n743) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n741), .ZN(n742) );
  NOR2_X1 U823 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U824 ( .A1(n745), .A2(n522), .ZN(n746) );
  NAND2_X1 U825 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U826 ( .A(n747), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U827 ( .A1(G8), .A2(n748), .ZN(n753) );
  INV_X1 U828 ( .A(n749), .ZN(n750) );
  NOR2_X1 U829 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U830 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U831 ( .A1(n755), .A2(n754), .ZN(n764) );
  NOR2_X1 U832 ( .A1(G303), .A2(G2090), .ZN(n756) );
  NAND2_X1 U833 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U834 ( .A(n757), .B(KEYINPUT98), .ZN(n758) );
  NAND2_X1 U835 ( .A1(n764), .A2(n758), .ZN(n759) );
  NAND2_X1 U836 ( .A1(n759), .A2(n777), .ZN(n773) );
  NOR2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n1012) );
  NOR2_X1 U838 ( .A1(G303), .A2(G1971), .ZN(n760) );
  NOR2_X1 U839 ( .A1(n1012), .A2(n760), .ZN(n762) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n761) );
  AND2_X1 U841 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U842 ( .A1(n764), .A2(n763), .ZN(n771) );
  NAND2_X1 U843 ( .A1(G288), .A2(G1976), .ZN(n1014) );
  INV_X1 U844 ( .A(n1014), .ZN(n765) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n520), .ZN(n767) );
  NAND2_X1 U846 ( .A1(n1012), .A2(KEYINPUT33), .ZN(n766) );
  OR2_X1 U847 ( .A1(n767), .A2(n523), .ZN(n769) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n1004) );
  INV_X1 U849 ( .A(n1004), .ZN(n768) );
  NOR2_X1 U850 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U851 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U852 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U854 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  XNOR2_X1 U855 ( .A(KEYINPUT100), .B(n779), .ZN(n813) );
  NAND2_X1 U856 ( .A1(G117), .A2(n898), .ZN(n786) );
  NAND2_X1 U857 ( .A1(G129), .A2(n873), .ZN(n781) );
  NAND2_X1 U858 ( .A1(G141), .A2(n621), .ZN(n780) );
  NAND2_X1 U859 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U860 ( .A1(n894), .A2(G105), .ZN(n782) );
  XOR2_X1 U861 ( .A(KEYINPUT38), .B(n782), .Z(n783) );
  NOR2_X1 U862 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U863 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U864 ( .A(n787), .B(KEYINPUT84), .ZN(n889) );
  NAND2_X1 U865 ( .A1(G1996), .A2(n889), .ZN(n796) );
  NAND2_X1 U866 ( .A1(G119), .A2(n873), .ZN(n789) );
  NAND2_X1 U867 ( .A1(G131), .A2(n621), .ZN(n788) );
  NAND2_X1 U868 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U869 ( .A1(G107), .A2(n898), .ZN(n790) );
  XNOR2_X1 U870 ( .A(KEYINPUT83), .B(n790), .ZN(n791) );
  NOR2_X1 U871 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U872 ( .A1(n894), .A2(G95), .ZN(n793) );
  NAND2_X1 U873 ( .A1(n794), .A2(n793), .ZN(n888) );
  NAND2_X1 U874 ( .A1(G1991), .A2(n888), .ZN(n795) );
  NAND2_X1 U875 ( .A1(n796), .A2(n795), .ZN(n975) );
  NOR2_X1 U876 ( .A1(n798), .A2(n797), .ZN(n827) );
  NAND2_X1 U877 ( .A1(n975), .A2(n827), .ZN(n799) );
  XNOR2_X1 U878 ( .A(n799), .B(KEYINPUT85), .ZN(n819) );
  XOR2_X1 U879 ( .A(KEYINPUT86), .B(n819), .Z(n810) );
  XNOR2_X1 U880 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NAND2_X1 U881 ( .A1(G104), .A2(n894), .ZN(n801) );
  NAND2_X1 U882 ( .A1(G140), .A2(n621), .ZN(n800) );
  NAND2_X1 U883 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n802), .ZN(n808) );
  NAND2_X1 U885 ( .A1(G128), .A2(n616), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G116), .A2(n898), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U888 ( .A(KEYINPUT35), .B(n805), .Z(n806) );
  XNOR2_X1 U889 ( .A(KEYINPUT82), .B(n806), .ZN(n807) );
  NOR2_X1 U890 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n809), .ZN(n906) );
  NOR2_X1 U892 ( .A1(n825), .A2(n906), .ZN(n994) );
  NAND2_X1 U893 ( .A1(n827), .A2(n994), .ZN(n822) );
  NAND2_X1 U894 ( .A1(n810), .A2(n822), .ZN(n811) );
  XOR2_X1 U895 ( .A(KEYINPUT87), .B(n811), .Z(n812) );
  NOR2_X1 U896 ( .A1(n813), .A2(n812), .ZN(n815) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n1009) );
  NAND2_X1 U898 ( .A1(n1009), .A2(n827), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n815), .A2(n814), .ZN(n830) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n889), .ZN(n984) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n888), .ZN(n976) );
  NOR2_X1 U903 ( .A1(n816), .A2(n976), .ZN(n817) );
  XOR2_X1 U904 ( .A(KEYINPUT101), .B(n817), .Z(n818) );
  NOR2_X1 U905 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U906 ( .A1(n984), .A2(n820), .ZN(n821) );
  XNOR2_X1 U907 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U908 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U909 ( .A(n824), .B(KEYINPUT102), .ZN(n826) );
  NAND2_X1 U910 ( .A1(n825), .A2(n906), .ZN(n991) );
  NAND2_X1 U911 ( .A1(n826), .A2(n991), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U913 ( .A1(n830), .A2(n829), .ZN(n832) );
  XOR2_X1 U914 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n831) );
  XNOR2_X1 U915 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U918 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U920 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n839), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2096), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U929 ( .A(G2090), .B(G2678), .ZN(n840) );
  XNOR2_X1 U930 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U931 ( .A(n842), .B(KEYINPUT104), .Z(n844) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U933 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U934 ( .A(KEYINPUT42), .B(G2100), .Z(n846) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n845) );
  XNOR2_X1 U936 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U937 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U938 ( .A(G1971), .B(G1956), .Z(n850) );
  XNOR2_X1 U939 ( .A(G1991), .B(G1966), .ZN(n849) );
  XNOR2_X1 U940 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U941 ( .A(G1976), .B(G1961), .Z(n852) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1981), .ZN(n851) );
  XNOR2_X1 U943 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U944 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U946 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U947 ( .A(G1996), .B(G2474), .Z(n857) );
  XNOR2_X1 U948 ( .A(n858), .B(n857), .ZN(G229) );
  XNOR2_X1 U949 ( .A(G286), .B(n1019), .ZN(n860) );
  XNOR2_X1 U950 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U951 ( .A(n1007), .B(G171), .Z(n861) );
  XNOR2_X1 U952 ( .A(n862), .B(n861), .ZN(n863) );
  NOR2_X1 U953 ( .A1(G37), .A2(n863), .ZN(n864) );
  XOR2_X1 U954 ( .A(KEYINPUT113), .B(n864), .Z(G397) );
  NAND2_X1 U955 ( .A1(G112), .A2(n898), .ZN(n865) );
  XNOR2_X1 U956 ( .A(n865), .B(KEYINPUT106), .ZN(n868) );
  NAND2_X1 U957 ( .A1(G124), .A2(n873), .ZN(n866) );
  XNOR2_X1 U958 ( .A(n866), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U959 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U960 ( .A1(G100), .A2(n894), .ZN(n870) );
  NAND2_X1 U961 ( .A1(G136), .A2(n621), .ZN(n869) );
  NAND2_X1 U962 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U963 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G130), .A2(n873), .ZN(n875) );
  NAND2_X1 U965 ( .A1(G118), .A2(n898), .ZN(n874) );
  NAND2_X1 U966 ( .A1(n875), .A2(n874), .ZN(n882) );
  XNOR2_X1 U967 ( .A(KEYINPUT108), .B(KEYINPUT45), .ZN(n880) );
  NAND2_X1 U968 ( .A1(n621), .A2(G142), .ZN(n878) );
  NAND2_X1 U969 ( .A1(n894), .A2(G106), .ZN(n876) );
  XOR2_X1 U970 ( .A(KEYINPUT107), .B(n876), .Z(n877) );
  NAND2_X1 U971 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U972 ( .A(n880), .B(n879), .Z(n881) );
  NOR2_X1 U973 ( .A1(n882), .A2(n881), .ZN(n886) );
  XOR2_X1 U974 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n884) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n883) );
  XNOR2_X1 U976 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U977 ( .A(n886), .B(n885), .Z(n887) );
  XNOR2_X1 U978 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U979 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U980 ( .A(G160), .B(G164), .ZN(n891) );
  XNOR2_X1 U981 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U982 ( .A(n893), .B(n974), .Z(n905) );
  NAND2_X1 U983 ( .A1(G103), .A2(n894), .ZN(n896) );
  NAND2_X1 U984 ( .A1(G139), .A2(n621), .ZN(n895) );
  NAND2_X1 U985 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U986 ( .A(KEYINPUT109), .B(n897), .Z(n903) );
  NAND2_X1 U987 ( .A1(G127), .A2(n873), .ZN(n900) );
  NAND2_X1 U988 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U989 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U991 ( .A1(n903), .A2(n902), .ZN(n979) );
  XNOR2_X1 U992 ( .A(G162), .B(n979), .ZN(n904) );
  XNOR2_X1 U993 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U994 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U995 ( .A1(G37), .A2(n908), .ZN(n909) );
  XNOR2_X1 U996 ( .A(KEYINPUT112), .B(n909), .ZN(G395) );
  XOR2_X1 U997 ( .A(G2451), .B(G2430), .Z(n911) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2443), .ZN(n910) );
  XNOR2_X1 U999 ( .A(n911), .B(n910), .ZN(n917) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n913) );
  XNOR2_X1 U1001 ( .A(G1348), .B(G1341), .ZN(n912) );
  XNOR2_X1 U1002 ( .A(n913), .B(n912), .ZN(n915) );
  XOR2_X1 U1003 ( .A(G2446), .B(G2427), .Z(n914) );
  XNOR2_X1 U1004 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1005 ( .A(n917), .B(n916), .Z(n918) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n918), .ZN(n924) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1010 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1011 ( .A1(G397), .A2(G395), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n924), .ZN(G401) );
  INV_X1 U1016 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G21), .ZN(n926) );
  XNOR2_X1 U1018 ( .A(G1961), .B(G5), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n936) );
  XOR2_X1 U1020 ( .A(G1348), .B(KEYINPUT59), .Z(n927) );
  XNOR2_X1 U1021 ( .A(G4), .B(n927), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(G20), .B(G1956), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(G1981), .B(G6), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(G19), .B(G1341), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1028 ( .A(KEYINPUT60), .B(n934), .Z(n935) );
  NAND2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n943) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(G23), .B(G1976), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n941), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT61), .B(n944), .Z(n945) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n945), .ZN(n946) );
  XOR2_X1 U1039 ( .A(KEYINPUT127), .B(n946), .Z(n1002) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n961) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT116), .B(n949), .ZN(n956) );
  XOR2_X1 U1045 ( .A(G1991), .B(G25), .Z(n950) );
  NAND2_X1 U1046 ( .A1(n950), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G27), .B(n951), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT117), .B(n952), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G32), .B(G1996), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n959), .B(KEYINPUT53), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(n967) );
  XOR2_X1 U1055 ( .A(G2090), .B(G35), .Z(n965) );
  XOR2_X1 U1056 ( .A(G2084), .B(KEYINPUT120), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G34), .B(n962), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT54), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n968), .ZN(n970) );
  INV_X1 U1062 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n971), .A2(G11), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT121), .ZN(n1000) );
  XNOR2_X1 U1066 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n996) );
  XOR2_X1 U1067 ( .A(G2084), .B(G160), .Z(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n990) );
  XOR2_X1 U1071 ( .A(G2072), .B(n979), .Z(n981) );
  XOR2_X1 U1072 ( .A(G164), .B(G2078), .Z(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT50), .B(n982), .ZN(n988) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT51), .B(n985), .Z(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT114), .B(n986), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n996), .B(n995), .ZN(n997) );
  OR2_X1 U1084 ( .A1(KEYINPUT55), .A2(n997), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(G29), .A2(n998), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1032) );
  XNOR2_X1 U1088 ( .A(G16), .B(KEYINPUT56), .ZN(n1029) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(KEYINPUT122), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1006), .B(KEYINPUT57), .ZN(n1027) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G166), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1025) );
  XOR2_X1 U1097 ( .A(n1012), .B(KEYINPUT124), .Z(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1015), .B(KEYINPUT125), .ZN(n1023) );
  XNOR2_X1 U1100 ( .A(G171), .B(G1961), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G1956), .B(KEYINPUT123), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1016), .B(G299), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(G1341), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1108 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1109 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1110 ( .A(n1030), .B(KEYINPUT126), .ZN(n1031) );
  NAND2_X1 U1111 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

