//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(new_n203), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT93), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(G1gat), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(new_n221), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(new_n217), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT93), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n214), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n219), .A2(new_n227), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n202), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n228), .B(new_n227), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n232), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n230), .A2(new_n228), .ZN(new_n238));
  INV_X1    g037(.A(new_n227), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n218), .B2(KEYINPUT93), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT18), .B(new_n232), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n241), .A3(new_n248), .A4(new_n237), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT94), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G64gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G71gat), .B(G78gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G127gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n227), .B1(new_n260), .B2(new_n261), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G183gat), .B(G211gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT95), .B(G155gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n265), .A2(new_n268), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n271));
  NAND2_X1  g070(.A1(G231gat), .A2(G233gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OR3_X1    g073(.A1(new_n269), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n269), .B2(new_n270), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT97), .B(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT98), .B(G92gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT7), .ZN(new_n282));
  INV_X1    g081(.A(G99gat), .ZN(new_n283));
  INV_X1    g082(.A(G106gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT8), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G99gat), .B(G106gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT17), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(new_n228), .ZN(new_n290));
  XOR2_X1   g089(.A(G190gat), .B(G218gat), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT41), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OR3_X1    g095(.A1(new_n290), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n290), .B2(new_n296), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT96), .B(G134gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n295), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n290), .A2(new_n292), .A3(new_n296), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(KEYINPUT99), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n299), .B(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n277), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G120gat), .B(G148gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G204gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G230gat), .ZN(new_n314));
  INV_X1    g113(.A(G233gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n286), .B(new_n287), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n260), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n288), .A2(new_n259), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT10), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n322), .A3(new_n320), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n288), .A2(KEYINPUT10), .A3(new_n259), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT100), .B1(new_n325), .B2(new_n317), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT100), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n327), .B(new_n316), .C1(new_n323), .C2(new_n324), .ZN(new_n328));
  OAI221_X1 g127(.A(new_n313), .B1(new_n317), .B2(new_n321), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n323), .A2(new_n324), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n316), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n321), .A2(new_n317), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n312), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(new_n333), .A3(KEYINPUT101), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n333), .A2(KEYINPUT101), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n307), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  NAND3_X1  g137(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(G183gat), .B2(G190gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT64), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  OR2_X1    g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n339), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT23), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(KEYINPUT23), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n338), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT67), .ZN(new_n356));
  INV_X1    g155(.A(new_n340), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n338), .B1(new_n360), .B2(KEYINPUT69), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n357), .B(new_n362), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(new_n354), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n338), .C1(new_n347), .C2(new_n354), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n356), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(G127gat), .A2(G134gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(G127gat), .A2(G134gat), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n369), .A2(KEYINPUT70), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT70), .B1(new_n369), .B2(new_n370), .ZN(new_n372));
  INV_X1    g171(.A(G120gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(G113gat), .ZN(new_n374));
  INV_X1    g173(.A(G113gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(G120gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n371), .A2(new_n372), .B1(new_n377), .B2(KEYINPUT1), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT1), .B1(new_n369), .B2(new_n370), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n375), .B2(G120gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n383), .B2(new_n374), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n386));
  OR3_X1    g185(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n350), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT27), .B(G183gat), .ZN(new_n390));
  INV_X1    g189(.A(G190gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT28), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT28), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n388), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n368), .A2(new_n385), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n385), .B1(new_n368), .B2(new_n395), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G227gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(new_n315), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT34), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT34), .ZN(new_n402));
  INV_X1    g201(.A(new_n400), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n403), .C1(new_n396), .C2(new_n397), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(G71gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(new_n283), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n368), .A2(new_n395), .ZN(new_n410));
  INV_X1    g209(.A(new_n385), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n368), .A2(new_n385), .A3(new_n395), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n400), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT72), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT72), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n412), .A2(new_n416), .A3(new_n400), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT32), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT33), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n409), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n408), .A2(KEYINPUT33), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n419), .B(new_n423), .C1(new_n415), .C2(new_n417), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n405), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n416), .B1(new_n398), .B2(new_n400), .ZN(new_n426));
  INV_X1    g225(.A(new_n417), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n408), .ZN(new_n429));
  INV_X1    g228(.A(new_n405), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n418), .A2(KEYINPUT32), .A3(new_n422), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n432), .A3(KEYINPUT73), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n429), .B2(new_n431), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT36), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n425), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G226gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n410), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT29), .B1(new_n368), .B2(new_n395), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n443), .B(KEYINPUT77), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n410), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n441), .ZN(new_n449));
  XNOR2_X1  g248(.A(G211gat), .B(G218gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(G197gat), .B(G204gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT22), .ZN(new_n452));
  INV_X1    g251(.A(G211gat), .ZN(new_n453));
  INV_X1    g252(.A(G218gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT75), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n450), .B(KEYINPUT74), .Z(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n449), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT76), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n410), .A2(new_n463), .A3(new_n442), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n447), .B2(new_n441), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(new_n443), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n467), .B2(new_n461), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT30), .ZN(new_n469));
  XOR2_X1   g268(.A(G8gat), .B(G36gat), .Z(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(G64gat), .ZN(new_n471));
  INV_X1    g270(.A(G92gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n445), .A2(new_n461), .A3(new_n449), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n443), .B(KEYINPUT76), .C1(new_n442), .C2(new_n444), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n461), .B1(new_n477), .B2(new_n464), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n462), .B(new_n473), .C1(new_n467), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT2), .ZN(new_n484));
  INV_X1    g283(.A(G148gat), .ZN(new_n485));
  OR2_X1    g284(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(G141gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT81), .B(new_n484), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G141gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G148gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT79), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT2), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n483), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(G155gat), .A2(G162gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(G155gat), .A2(G162gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n495), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT78), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT81), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n484), .C1(new_n488), .C2(new_n490), .ZN(new_n509));
  INV_X1    g308(.A(new_n503), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n411), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n385), .A3(new_n511), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n482), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT83), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n518));
  INV_X1    g317(.A(new_n482), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n507), .A2(new_n385), .A3(new_n511), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n385), .B1(new_n507), .B2(new_n511), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT5), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT4), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n521), .A2(new_n526), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT3), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n385), .B1(new_n512), .B2(new_n529), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n527), .A2(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(new_n519), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n525), .A2(KEYINPUT5), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n517), .A2(KEYINPUT82), .A3(new_n524), .ZN(new_n536));
  OAI221_X1 g335(.A(new_n482), .B1(new_n531), .B2(new_n532), .C1(new_n527), .C2(new_n528), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G1gat), .B(G29gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT0), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G57gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(G85gat), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT6), .ZN(new_n545));
  INV_X1    g344(.A(new_n543), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n535), .A2(new_n546), .A3(new_n538), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n535), .A2(new_n538), .A3(KEYINPUT6), .A4(new_n546), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n475), .A2(new_n481), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G22gat), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n507), .A2(new_n511), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT29), .B1(new_n457), .B2(new_n460), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(KEYINPUT3), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT85), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n461), .B1(new_n530), .B2(new_n446), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G228gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(new_n315), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT85), .B(new_n552), .C1(new_n553), .C2(KEYINPUT3), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n556), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n459), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n457), .B1(new_n450), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n446), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n512), .B1(new_n565), .B2(new_n529), .ZN(new_n566));
  OAI22_X1  g365(.A1(new_n566), .A2(new_n557), .B1(new_n559), .B2(new_n315), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n551), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n567), .A3(new_n551), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G78gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G50gat), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n569), .A2(new_n576), .A3(new_n570), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n550), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT87), .B1(new_n440), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n548), .A2(new_n549), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n476), .B2(new_n478), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT90), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n468), .A2(new_n589), .A3(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n461), .B1(new_n445), .B2(new_n449), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n592), .B1(new_n461), .B2(new_n467), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT38), .B1(new_n593), .B2(KEYINPUT37), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n473), .A3(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n476), .A2(new_n478), .A3(new_n586), .ZN(new_n596));
  AOI211_X1 g395(.A(new_n474), .B(new_n596), .C1(new_n588), .C2(new_n590), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT38), .B1(new_n468), .B2(new_n474), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n585), .B(new_n595), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n533), .A2(new_n519), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n513), .A2(new_n482), .A3(new_n514), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT39), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT88), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT88), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT39), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n533), .A2(new_n607), .A3(new_n519), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n606), .A2(KEYINPUT40), .A3(new_n543), .A4(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT89), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n543), .A3(new_n608), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n614), .A2(new_n547), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n481), .A2(new_n475), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n580), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n584), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n580), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n437), .A4(new_n439), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n583), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n421), .A2(new_n424), .A3(new_n405), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n434), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n425), .A2(new_n432), .A3(KEYINPUT91), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n628), .A2(new_n550), .A3(new_n581), .A4(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT35), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n621), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n580), .B1(new_n433), .B2(new_n436), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n254), .B(new_n337), .C1(new_n625), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n585), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G1gat), .ZN(G1324gat));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n254), .B1(new_n625), .B2(new_n634), .ZN(new_n639));
  INV_X1    g438(.A(new_n337), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n618), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(new_n643), .A3(new_n618), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n222), .A2(KEYINPUT42), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT16), .B(G8gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT103), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n635), .A2(KEYINPUT42), .A3(new_n618), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n638), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n652), .A2(new_n649), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(KEYINPUT104), .A3(new_n646), .A4(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n628), .A2(new_n629), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(G15gat), .B1(new_n635), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n440), .A2(G15gat), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n635), .B2(new_n661), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n625), .A2(new_n634), .ZN(new_n663));
  INV_X1    g462(.A(new_n254), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n580), .A4(new_n640), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT105), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n639), .A2(new_n668), .A3(new_n580), .A4(new_n640), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n667), .B1(new_n666), .B2(new_n669), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n671), .A2(new_n672), .A3(new_n551), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n666), .A2(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT43), .ZN(new_n675));
  AOI21_X1  g474(.A(G22gat), .B1(new_n675), .B2(new_n670), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n673), .A2(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n277), .ZN(new_n678));
  INV_X1    g477(.A(new_n336), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n639), .A2(new_n306), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n207), .A3(new_n585), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  INV_X1    g482(.A(new_n440), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n550), .B2(new_n581), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n621), .A2(KEYINPUT106), .A3(new_n580), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n620), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n634), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n690), .B2(new_n306), .ZN(new_n691));
  INV_X1    g490(.A(new_n306), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n625), .B2(new_n634), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n252), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT107), .B1(new_n700), .B2(new_n584), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n697), .A2(new_n702), .A3(new_n585), .A4(new_n699), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(G29gat), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n704), .ZN(G1328gat));
  AND3_X1   g504(.A1(new_n681), .A2(new_n208), .A3(new_n618), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n700), .B2(new_n617), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n707), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  NAND4_X1  g510(.A1(new_n697), .A2(G43gat), .A3(new_n440), .A4(new_n699), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n639), .A2(new_n659), .A3(new_n306), .A4(new_n680), .ZN(new_n713));
  INV_X1    g512(.A(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n713), .A2(new_n714), .B1(new_n715), .B2(KEYINPUT47), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(KEYINPUT47), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT109), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n717), .B(new_n719), .ZN(G1330gat));
  NOR2_X1   g519(.A1(new_n581), .A2(G50gat), .ZN(new_n721));
  AND4_X1   g520(.A1(new_n639), .A2(new_n306), .A3(new_n680), .A4(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR4_X1   g522(.A1(new_n691), .A2(new_n696), .A3(new_n581), .A4(new_n698), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n630), .A2(new_n631), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n632), .A2(new_n633), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n440), .B1(new_n686), .B2(new_n687), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n620), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n693), .B1(new_n733), .B2(new_n692), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n663), .A2(new_n694), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n734), .A2(new_n580), .A3(new_n735), .A4(new_n699), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n722), .B1(new_n736), .B2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n737), .A2(KEYINPUT110), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n728), .A2(new_n739), .ZN(G1331gat));
  INV_X1    g539(.A(new_n252), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n690), .A2(new_n741), .A3(new_n307), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n679), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n585), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n617), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n744), .A2(G71gat), .A3(new_n440), .ZN(new_n752));
  INV_X1    g551(.A(G71gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n743), .B2(new_n658), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT50), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n752), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1334gat));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n581), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT111), .B(G78gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1335gat));
  AOI21_X1  g561(.A(new_n692), .B1(new_n689), .B2(new_n634), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n678), .A2(new_n252), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n763), .A2(KEYINPUT51), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT51), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n585), .A3(new_n278), .A4(new_n679), .ZN(new_n769));
  INV_X1    g568(.A(new_n764), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n691), .A2(new_n696), .A3(new_n336), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(KEYINPUT112), .A3(new_n585), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n734), .A2(new_n679), .A3(new_n735), .A4(new_n764), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n584), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(new_n776), .B2(new_n278), .ZN(G1336gat));
  AOI21_X1  g576(.A(new_n279), .B1(new_n771), .B2(new_n618), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n617), .A2(G92gat), .A3(new_n336), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT113), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT52), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n279), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n774), .B2(new_n617), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n784), .B(new_n785), .C1(new_n767), .C2(new_n780), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n774), .B2(new_n684), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n768), .A2(new_n283), .A3(new_n659), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n336), .ZN(G1338gat));
  XOR2_X1   g589(.A(KEYINPUT114), .B(G106gat), .Z(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n771), .B2(new_n580), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n581), .A2(G106gat), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n679), .B(new_n794), .C1(new_n765), .C2(new_n766), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n774), .B2(new_n581), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n796), .A3(new_n800), .A4(new_n795), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1339gat));
  NAND2_X1  g601(.A1(new_n330), .A2(new_n316), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT54), .B(new_n803), .C1(new_n326), .C2(new_n328), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n313), .B1(new_n331), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n804), .B2(new_n806), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n252), .B(new_n329), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n235), .A2(new_n236), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n238), .A2(new_n240), .A3(new_n232), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n247), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n251), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n334), .A2(new_n335), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n306), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n329), .B(new_n814), .C1(new_n808), .C2(new_n809), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n692), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n277), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n307), .A2(new_n741), .A3(new_n336), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n658), .A2(new_n580), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n618), .A2(new_n584), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n254), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n580), .B1(new_n819), .B2(new_n820), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n433), .A2(new_n436), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n823), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n252), .A2(new_n375), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT116), .Z(new_n831));
  OAI21_X1  g630(.A(new_n825), .B1(new_n829), .B2(new_n831), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n824), .B2(new_n336), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n679), .A2(new_n373), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n829), .B2(new_n834), .ZN(G1341gat));
  INV_X1    g634(.A(new_n829), .ZN(new_n836));
  AOI21_X1  g635(.A(G127gat), .B1(new_n836), .B2(new_n678), .ZN(new_n837));
  INV_X1    g636(.A(new_n824), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(G127gat), .A3(new_n678), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(G1342gat));
  OR3_X1    g641(.A1(new_n829), .A2(G134gat), .A3(new_n692), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n824), .B2(new_n692), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n843), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n844), .B(new_n845), .C1(new_n848), .C2(new_n849), .ZN(G1343gat));
  AND2_X1   g649(.A1(new_n486), .A2(new_n487), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n684), .A2(new_n585), .A3(new_n617), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n329), .B1(new_n808), .B2(new_n809), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n815), .B1(new_n254), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n692), .ZN(new_n858));
  INV_X1    g657(.A(new_n818), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n678), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n820), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n580), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n821), .A2(new_n580), .ZN(new_n863));
  XOR2_X1   g662(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n855), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n851), .B1(new_n868), .B2(new_n254), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n581), .B1(new_n819), .B2(new_n820), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n585), .A3(new_n684), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n618), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n492), .A3(new_n664), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n869), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n867), .A2(new_n252), .A3(new_n854), .A4(new_n853), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n879), .A2(new_n880), .A3(new_n851), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n879), .B2(new_n851), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n871), .A2(G141gat), .A3(new_n254), .A4(new_n618), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n878), .B1(new_n884), .B2(new_n877), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n875), .A2(new_n485), .A3(new_n679), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n855), .A2(new_n867), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n485), .C1(new_n887), .C2(new_n679), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n864), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n818), .B1(new_n857), .B2(new_n692), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n891), .A2(new_n678), .B1(new_n664), .B2(new_n337), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n580), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n679), .A3(new_n855), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n889), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n886), .B1(new_n888), .B2(new_n896), .ZN(G1345gat));
  AND3_X1   g696(.A1(new_n887), .A2(G155gat), .A3(new_n678), .ZN(new_n898));
  AOI21_X1  g697(.A(G155gat), .B1(new_n875), .B2(new_n678), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT123), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n887), .A2(G155gat), .A3(new_n678), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n875), .A2(new_n678), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(G155gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n904), .ZN(G1346gat));
  AND3_X1   g704(.A1(new_n887), .A2(G162gat), .A3(new_n306), .ZN(new_n906));
  AOI21_X1  g705(.A(G162gat), .B1(new_n875), .B2(new_n306), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1347gat));
  NOR3_X1   g707(.A1(new_n658), .A2(new_n585), .A3(new_n617), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT124), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(KEYINPUT124), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n826), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n254), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n585), .A2(new_n617), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n828), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n741), .A2(G169gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1348gat));
  NOR3_X1   g716(.A1(new_n912), .A2(new_n309), .A3(new_n336), .ZN(new_n918));
  INV_X1    g717(.A(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n679), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n920), .B2(new_n309), .ZN(G1349gat));
  OAI21_X1  g720(.A(G183gat), .B1(new_n912), .B2(new_n277), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n678), .A2(new_n390), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n391), .A3(new_n306), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n306), .A3(new_n826), .A4(new_n911), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(G190gat), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n928), .A2(new_n927), .A3(G190gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT125), .Z(G1351gat));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n890), .B(new_n933), .C1(new_n893), .C2(KEYINPUT57), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n892), .B2(new_n580), .ZN(new_n935));
  INV_X1    g734(.A(new_n890), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT126), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n684), .A2(new_n914), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n664), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G197gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n863), .A2(new_n939), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n944), .A3(new_n252), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(G1352gat));
  NAND4_X1  g745(.A1(new_n938), .A2(KEYINPUT127), .A3(new_n679), .A4(new_n940), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n934), .A2(new_n937), .A3(new_n679), .A4(new_n940), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n947), .A2(G204gat), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n943), .A2(new_n311), .A3(new_n679), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n943), .A2(new_n453), .A3(new_n678), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n894), .A2(new_n678), .A3(new_n940), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n943), .B2(new_n306), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n938), .A2(new_n940), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n692), .A2(new_n454), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1355gat));
endmodule


