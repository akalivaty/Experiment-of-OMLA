//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(KEYINPUT76), .A3(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n211), .A2(new_n213), .B1(KEYINPUT2), .B2(new_n205), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n207), .B(new_n206), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G113gat), .B(G120gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g022(.A(G127gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225));
  INV_X1    g024(.A(G134gat), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G120gat), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n225), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n223), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n224), .B1(new_n223), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n219), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT78), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n236), .B(new_n219), .C1(new_n232), .C2(new_n233), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n233), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n231), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n219), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n219), .A2(new_n244), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n238), .A2(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n247), .B2(new_n245), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT4), .B1(new_n235), .B2(new_n237), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n242), .B1(new_n241), .B2(new_n219), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n232), .A2(new_n233), .ZN(new_n257));
  INV_X1    g056(.A(new_n219), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n235), .A2(new_n237), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n249), .B1(new_n260), .B2(new_n252), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n256), .B1(new_n261), .B2(KEYINPUT79), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n251), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G85gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT81), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n268), .B(new_n251), .C1(new_n262), .C2(new_n263), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT81), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(new_n275), .A3(new_n269), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n269), .ZN(new_n278));
  XNOR2_X1  g077(.A(G197gat), .B(G204gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n281));
  INV_X1    g080(.A(G211gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n279), .B1(new_n285), .B2(KEYINPUT22), .ZN(new_n286));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n279), .B(new_n287), .C1(new_n285), .C2(KEYINPUT22), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G226gat), .ZN(new_n292));
  INV_X1    g091(.A(G233gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n298), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT27), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT28), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n311), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n318));
  NOR3_X1   g117(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n302), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT25), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n321), .A2(new_n302), .A3(new_n323), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n318), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n310), .A3(KEYINPUT65), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n332), .A3(new_n316), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n326), .B(new_n327), .C1(new_n329), .C2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n314), .A2(new_n325), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n318), .B(KEYINPUT64), .ZN(new_n337));
  INV_X1    g136(.A(new_n333), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n340));
  INV_X1    g139(.A(new_n318), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n306), .A3(new_n310), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n341), .A2(new_n343), .A3(new_n315), .A4(new_n316), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n339), .A2(new_n340), .B1(new_n345), .B2(KEYINPUT25), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n314), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n295), .B1(new_n336), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n294), .A2(KEYINPUT29), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n314), .A2(new_n334), .A3(KEYINPUT72), .A4(new_n325), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n291), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n348), .A3(new_n350), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n294), .A3(new_n354), .ZN(new_n358));
  INV_X1    g157(.A(new_n291), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT74), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(new_n360), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(KEYINPUT37), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n369));
  NAND3_X1  g168(.A1(new_n357), .A2(new_n358), .A3(new_n291), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT37), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n347), .B1(new_n346), .B2(new_n314), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n294), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT72), .B1(new_n346), .B2(new_n314), .ZN(new_n375));
  INV_X1    g174(.A(new_n354), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n350), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n291), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n369), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n365), .B1(new_n368), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n356), .A2(new_n381), .A3(new_n360), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(new_n356), .B2(new_n360), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT37), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n368), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n369), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n380), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n277), .A2(new_n278), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n356), .A2(KEYINPUT30), .A3(new_n360), .A4(new_n364), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT75), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n359), .B1(new_n374), .B2(new_n377), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n356), .A2(new_n381), .A3(new_n360), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n397), .B2(new_n366), .ZN(new_n398));
  INV_X1    g197(.A(new_n365), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n248), .A2(new_n250), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT39), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n269), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n260), .A2(new_n252), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(KEYINPUT39), .C1(new_n248), .C2(new_n250), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n403), .A2(KEYINPUT40), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT40), .B1(new_n403), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n400), .A2(new_n408), .A3(new_n271), .A4(new_n276), .ZN(new_n409));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT80), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n410), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n219), .B2(new_n244), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n415), .A2(new_n291), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n289), .B2(new_n290), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n258), .B1(new_n417), .B2(KEYINPUT3), .ZN(new_n418));
  INV_X1    g217(.A(G22gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(KEYINPUT80), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n415), .B2(new_n291), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423));
  INV_X1    g222(.A(new_n290), .ZN(new_n424));
  INV_X1    g223(.A(new_n284), .ZN(new_n425));
  NOR2_X1   g224(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n426));
  OAI21_X1  g225(.A(G218gat), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT22), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n287), .B1(new_n429), .B2(new_n279), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n219), .B1(new_n431), .B2(new_n244), .ZN(new_n432));
  OAI21_X1  g231(.A(G22gat), .B1(new_n422), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT31), .B(G50gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n421), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n421), .B2(new_n433), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n414), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n434), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n433), .A3(new_n435), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n413), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n389), .A2(new_n409), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G15gat), .B(G43gat), .Z(new_n445));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n257), .A2(new_n346), .A3(new_n314), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n335), .A2(new_n241), .ZN(new_n450));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n451), .B2(KEYINPUT69), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n449), .A2(new_n450), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  AOI211_X1 g259(.A(new_n452), .B(new_n457), .C1(new_n449), .C2(new_n450), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n455), .A2(new_n460), .A3(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(new_n453), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT32), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n460), .A2(new_n461), .ZN(new_n468));
  INV_X1    g267(.A(new_n455), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n467), .A2(KEYINPUT36), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT36), .B1(new_n467), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n390), .B(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n366), .B1(new_n382), .B2(new_n383), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT30), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n365), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n272), .A2(new_n273), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n256), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n268), .B1(new_n484), .B2(new_n251), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n278), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n438), .A2(new_n442), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n475), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n470), .A2(new_n471), .A3(new_n462), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n471), .B1(new_n470), .B2(new_n462), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n490), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n480), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n277), .A2(new_n278), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n443), .A2(new_n467), .A3(new_n472), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n400), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n444), .A2(new_n489), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G197gat), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT11), .B(G169gat), .Z(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(KEYINPUT12), .Z(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT13), .Z(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT84), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT84), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT85), .B(G29gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  INV_X1    g322(.A(G43gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(G50gat), .ZN(new_n525));
  INV_X1    g324(.A(G50gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(G43gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n514), .A2(new_n508), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n520), .A2(new_n517), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n532), .A2(G1gat), .ZN(new_n536));
  OAI21_X1  g335(.A(G8gat), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n538), .B(new_n539), .C1(G1gat), .C2(new_n532), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n522), .A2(new_n530), .B1(new_n537), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n507), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(KEYINPUT88), .B(new_n507), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n508), .A2(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n549), .A2(new_n511), .B1(G36gat), .B2(new_n516), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n530), .B(KEYINPUT17), .C1(new_n520), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n522), .A2(KEYINPUT87), .A3(KEYINPUT17), .A4(new_n530), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT86), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n520), .A2(new_n517), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n528), .A2(new_n529), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n557), .A2(new_n558), .B1(new_n518), .B2(new_n521), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n556), .B1(new_n559), .B2(KEYINPUT17), .ZN(new_n560));
  INV_X1    g359(.A(new_n541), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n531), .A2(KEYINPUT86), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n555), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n543), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n506), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n543), .B1(G229gat), .B2(G233gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT18), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n505), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n569), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n505), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n567), .A4(new_n548), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n576), .A3(KEYINPUT89), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT89), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n578), .B(new_n505), .C1(new_n568), .C2(new_n570), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n500), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n583));
  XOR2_X1   g382(.A(G99gat), .B(G106gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT8), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(G99gat), .B2(G106gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT94), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G99gat), .A2(G106gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT8), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  INV_X1    g392(.A(G92gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n585), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n584), .B(new_n602), .C1(new_n589), .C2(new_n596), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n555), .A2(new_n560), .A3(new_n563), .A4(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n606), .A2(new_n531), .B1(KEYINPUT41), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT95), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(new_n610), .A3(new_n613), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT96), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n615), .A2(KEYINPUT96), .A3(new_n619), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(new_n616), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G134gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n203), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n618), .A2(new_n624), .A3(new_n627), .A4(new_n620), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  OR2_X1    g431(.A1(G71gat), .A2(G78gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(G71gat), .A2(G78gat), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT9), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G57gat), .B(G64gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(KEYINPUT90), .ZN(new_n639));
  INV_X1    g438(.A(G57gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G64gat), .ZN(new_n641));
  INV_X1    g440(.A(G64gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(G57gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n643), .A3(KEYINPUT90), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n635), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n640), .A2(G64gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT91), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT91), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n641), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n634), .B1(new_n633), .B2(new_n636), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n561), .B1(new_n632), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT93), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n632), .ZN(new_n657));
  XNOR2_X1  g456(.A(G127gat), .B(G155gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n656), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT92), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n660), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n583), .B1(new_n631), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n629), .A2(new_n670), .A3(KEYINPUT98), .A4(new_n630), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n654), .B1(new_n604), .B2(new_n605), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT90), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n642), .A2(G57gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n647), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n644), .A3(new_n637), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n679), .A2(new_n635), .B1(new_n651), .B2(new_n652), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n592), .B1(new_n591), .B2(new_n595), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n603), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n584), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n597), .A2(new_n585), .A3(new_n603), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n674), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT99), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n674), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT10), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n675), .A2(new_n694), .A3(new_n686), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n680), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n687), .A2(KEYINPUT99), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n692), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n691), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n697), .B2(new_n687), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n672), .A2(new_n673), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n672), .A2(new_n707), .A3(new_n673), .A4(new_n704), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n582), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n486), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n400), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT101), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT101), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(G8gat), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT16), .B(G8gat), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n715), .B2(new_n716), .ZN(new_n721));
  OAI221_X1 g520(.A(new_n717), .B1(new_n714), .B2(new_n719), .C1(new_n721), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g521(.A(new_n710), .ZN(new_n723));
  INV_X1    g522(.A(new_n475), .ZN(new_n724));
  OAI21_X1  g523(.A(G15gat), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n490), .A2(new_n491), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(G15gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n723), .B2(new_n728), .ZN(G1326gat));
  NAND2_X1  g528(.A1(new_n710), .A2(new_n488), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT102), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT43), .B(G22gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1327gat));
  AND2_X1   g532(.A1(new_n629), .A2(new_n630), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n500), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n581), .A2(new_n670), .A3(new_n703), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n486), .A3(new_n516), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n444), .A2(new_n489), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n494), .A2(new_n499), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(KEYINPUT44), .A3(new_n631), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n500), .B2(new_n734), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n711), .A3(new_n736), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n516), .B1(new_n748), .B2(KEYINPUT103), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n740), .B(new_n753), .C1(new_n749), .C2(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1328gat));
  INV_X1    g554(.A(new_n737), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n513), .A3(new_n400), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT46), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n747), .A2(new_n736), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n513), .B1(new_n759), .B2(new_n400), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n758), .A2(new_n760), .ZN(G1329gat));
  NAND3_X1  g560(.A1(new_n759), .A2(G43gat), .A3(new_n475), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n524), .B1(new_n737), .B2(new_n727), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g564(.A1(new_n759), .A2(new_n488), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G50gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT48), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n756), .A2(new_n526), .A3(new_n488), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n767), .B(new_n770), .C1(new_n768), .C2(KEYINPUT48), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1331gat));
  AND2_X1   g573(.A1(new_n672), .A2(new_n673), .ZN(new_n775));
  AND4_X1   g574(.A1(new_n775), .A2(new_n743), .A3(new_n703), .A4(new_n581), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n711), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT106), .B(G57gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1332gat));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n400), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT49), .B(G64gat), .Z(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n780), .B2(new_n782), .ZN(G1333gat));
  NAND3_X1  g582(.A1(new_n776), .A2(G71gat), .A3(new_n475), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n776), .A2(new_n726), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  INV_X1    g585(.A(G71gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n785), .B2(KEYINPUT107), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n776), .A2(new_n488), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n580), .A2(new_n670), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n703), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT108), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n744), .A2(new_n746), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n744), .A2(new_n746), .A3(new_n798), .A4(new_n795), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n711), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n593), .B1(new_n800), .B2(KEYINPUT110), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(KEYINPUT110), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n735), .A2(new_n793), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n735), .A2(new_n805), .A3(new_n793), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n703), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n711), .A2(new_n593), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(G1336gat));
  INV_X1    g608(.A(new_n807), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n594), .A3(new_n400), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n797), .A2(new_n400), .A3(new_n799), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815));
  INV_X1    g614(.A(new_n796), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n594), .B1(new_n816), .B2(new_n400), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n811), .A2(new_n815), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n814), .A2(new_n815), .B1(new_n817), .B2(new_n818), .ZN(G1337gat));
  AND3_X1   g618(.A1(new_n797), .A2(new_n475), .A3(new_n799), .ZN(new_n820));
  XOR2_X1   g619(.A(KEYINPUT111), .B(G99gat), .Z(new_n821));
  NAND2_X1  g620(.A1(new_n726), .A2(new_n821), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n820), .A2(new_n821), .B1(new_n807), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT112), .ZN(G1338gat));
  NOR3_X1   g623(.A1(new_n807), .A2(G106gat), .A3(new_n443), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g625(.A(G106gat), .B1(new_n796), .B2(new_n443), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n797), .A2(new_n488), .A3(new_n799), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n829), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT113), .B1(new_n829), .B2(G106gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n831), .A3(new_n825), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(G1339gat));
  NAND2_X1  g633(.A1(new_n695), .A2(new_n696), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n674), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n695), .A2(new_n693), .A3(new_n696), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  XOR2_X1   g637(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n839));
  AOI21_X1  g638(.A(new_n691), .B1(new_n697), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n838), .A2(new_n840), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n838), .B2(new_n840), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n699), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n506), .B1(new_n564), .B2(new_n565), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n542), .A2(new_n543), .A3(new_n507), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n504), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n576), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n631), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n845), .A2(new_n579), .A3(new_n577), .A4(new_n847), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n703), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(KEYINPUT116), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n734), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT116), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT117), .B(new_n853), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n671), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n775), .A2(new_n704), .A3(new_n581), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n711), .A3(new_n492), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n486), .B1(new_n863), .B2(new_n864), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT119), .A3(new_n492), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n400), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n580), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n865), .B2(new_n443), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT118), .B(new_n488), .C1(new_n863), .C2(new_n864), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n486), .A2(new_n400), .A3(new_n727), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n581), .A2(new_n227), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n872), .B1(new_n879), .B2(new_n880), .ZN(G1340gat));
  AOI21_X1  g680(.A(G120gat), .B1(new_n871), .B2(new_n703), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n704), .A2(new_n229), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n879), .B2(new_n883), .ZN(G1341gat));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n870), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n670), .A3(new_n480), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT68), .B(G127gat), .Z(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n671), .A2(new_n887), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT120), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  INV_X1    g691(.A(new_n887), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n871), .B2(new_n670), .ZN(new_n894));
  NOR4_X1   g693(.A1(new_n876), .A2(new_n671), .A3(new_n878), .A4(new_n887), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(G1342gat));
  NAND2_X1  g696(.A1(new_n631), .A2(new_n480), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT121), .Z(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(G134gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n900), .A3(new_n902), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n631), .B(new_n877), .C1(new_n874), .C2(new_n875), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G134gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G134gat), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n904), .B(new_n905), .C1(new_n908), .C2(new_n909), .ZN(G1343gat));
  NAND3_X1  g709(.A1(new_n869), .A2(new_n488), .A3(new_n724), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n400), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n580), .A2(new_n210), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT124), .Z(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n475), .A2(new_n486), .A3(new_n400), .ZN(new_n916));
  INV_X1    g715(.A(new_n853), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n631), .B1(new_n854), .B2(new_n855), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n671), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n443), .B1(new_n864), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n443), .B1(new_n863), .B2(new_n864), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(new_n580), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n915), .B1(new_n925), .B2(new_n210), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT58), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(new_n915), .C1(new_n925), .C2(new_n210), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1344gat));
  NOR2_X1   g729(.A1(new_n704), .A2(G148gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n912), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n706), .A2(new_n708), .A3(new_n581), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n919), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n488), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n921), .ZN(new_n938));
  AOI211_X1 g737(.A(new_n921), .B(new_n443), .C1(new_n863), .C2(new_n864), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(KEYINPUT126), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n923), .A2(KEYINPUT126), .A3(KEYINPUT57), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n703), .B(new_n916), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n934), .B1(new_n942), .B2(G148gat), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT59), .B(new_n212), .C1(new_n924), .C2(new_n703), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n933), .B1(new_n943), .B2(new_n944), .ZN(G1345gat));
  NAND3_X1  g744(.A1(new_n912), .A2(new_n202), .A3(new_n670), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n924), .A2(new_n670), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(new_n202), .ZN(G1346gat));
  OR3_X1    g747(.A1(new_n911), .A2(G162gat), .A3(new_n899), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n924), .A2(new_n631), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n203), .ZN(G1347gat));
  AOI21_X1  g750(.A(new_n711), .B1(new_n863), .B2(new_n864), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n400), .A2(new_n492), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G169gat), .B1(new_n954), .B2(new_n580), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n711), .A2(new_n480), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n726), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n876), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n580), .A2(G169gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1348gat));
  INV_X1    g759(.A(G176gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n954), .A2(new_n961), .A3(new_n703), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n876), .A2(new_n704), .A3(new_n957), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n961), .ZN(G1349gat));
  AND3_X1   g763(.A1(new_n670), .A2(new_n307), .A3(new_n309), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n952), .A2(new_n953), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n957), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n670), .B(new_n969), .C1(new_n874), .C2(new_n875), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n970), .B2(G183gat), .ZN(new_n971));
  NOR2_X1   g770(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n310), .A3(new_n631), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n631), .B(new_n969), .C1(new_n874), .C2(new_n875), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n975), .A2(new_n976), .A3(G190gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n975), .B2(G190gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1351gat));
  NOR3_X1   g778(.A1(new_n475), .A2(new_n443), .A3(new_n480), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n952), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n580), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n940), .A2(new_n941), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n475), .A2(new_n711), .A3(new_n480), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n580), .A2(G197gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NAND3_X1  g786(.A1(new_n983), .A2(new_n703), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G204gat), .ZN(new_n989));
  INV_X1    g788(.A(G204gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n981), .A2(new_n990), .A3(new_n703), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  NAND2_X1  g791(.A1(new_n989), .A2(new_n992), .ZN(G1353gat));
  NAND4_X1  g792(.A1(new_n981), .A2(new_n670), .A3(new_n283), .A4(new_n284), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n670), .B(new_n984), .C1(new_n940), .C2(new_n941), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n631), .A3(new_n984), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G218gat), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n981), .A2(new_n280), .A3(new_n631), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


