//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1309, new_n1310, new_n1311, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  INV_X1    g0042(.A(G107), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G97), .ZN(new_n244));
  INV_X1    g0044(.A(G97), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G107), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n242), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n216), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n206), .B2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT8), .A2(G58), .ZN(new_n255));
  INV_X1    g0055(.A(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n255), .B1(new_n260), .B2(KEYINPUT8), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(new_n261), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT66), .B(G58), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n213), .B1(new_n266), .B2(new_n220), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n267), .A2(G20), .B1(G159), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT7), .B1(new_n272), .B2(new_n207), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(G68), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n269), .A2(new_n280), .A3(KEYINPUT16), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n252), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n276), .A2(new_n207), .A3(new_n277), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT7), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n278), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(KEYINPUT70), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G68), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT16), .B1(new_n289), .B2(new_n269), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n265), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n275), .A2(new_n222), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G223), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n276), .A2(new_n277), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT65), .B1(new_n298), .B2(new_n216), .ZN(new_n299));
  AND2_X1   g0099(.A1(G1), .A2(G13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT65), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT71), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n299), .A2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(G223), .ZN(new_n307));
  INV_X1    g0107(.A(G1698), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n294), .A2(G1698), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n309), .B(new_n310), .C1(new_n270), .C2(new_n271), .ZN(new_n311));
  INV_X1    g0111(.A(new_n292), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT71), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n306), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G274), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n300), .B2(new_n302), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n302), .A2(G1), .A3(G13), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G232), .A3(new_n318), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n305), .A2(new_n315), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n304), .B1(new_n312), .B2(new_n311), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n320), .A2(new_n322), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n291), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT18), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n291), .A2(new_n334), .A3(new_n331), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n282), .A2(new_n290), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n320), .A2(new_n322), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n305), .A2(new_n315), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n327), .B2(new_n328), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n336), .A2(KEYINPUT17), .A3(new_n265), .A4(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n265), .C1(new_n282), .C2(new_n290), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n333), .A2(new_n335), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n252), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n207), .A2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n261), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n264), .A2(new_n202), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n254), .B2(new_n202), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT9), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n296), .A2(G222), .A3(new_n308), .ZN(new_n358));
  INV_X1    g0158(.A(G77), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n296), .A2(G1698), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n358), .B1(new_n359), .B2(new_n296), .C1(new_n360), .C2(new_n307), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n306), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n321), .A2(new_n318), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT64), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT64), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n321), .A2(new_n365), .A3(new_n318), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G226), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n362), .A2(new_n320), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G200), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n356), .A2(KEYINPUT9), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n362), .A2(G190), .A3(new_n320), .A4(new_n368), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n357), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT10), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n370), .A4(new_n357), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n356), .B1(new_n369), .B2(new_n326), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G179), .B2(new_n369), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n253), .A2(G77), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G77), .B2(new_n263), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT8), .B(G58), .Z(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n349), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n252), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n367), .A2(G244), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n389), .A2(new_n320), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n296), .A2(G232), .A3(new_n308), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n391), .B1(new_n243), .B2(new_n296), .C1(new_n360), .C2(new_n221), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n306), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n390), .A2(G190), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n394), .B2(KEYINPUT67), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n340), .B1(new_n390), .B2(new_n393), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT67), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(new_n393), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n396), .A2(new_n397), .B1(new_n398), .B2(new_n337), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(new_n323), .A3(new_n393), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n387), .B1(new_n398), .B2(new_n326), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n395), .A2(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n378), .A2(new_n380), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n275), .A2(new_n245), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G226), .A2(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n232), .B2(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n406), .B2(new_n296), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n320), .B1(new_n407), .B2(new_n304), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n221), .B1(new_n364), .B2(new_n366), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT13), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n232), .A2(G1698), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(G226), .B2(G1698), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n413), .A2(new_n272), .B1(new_n275), .B2(new_n245), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n306), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n321), .A2(new_n365), .A3(new_n318), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n365), .B1(new_n321), .B2(new_n318), .ZN(new_n417));
  OAI21_X1  g0217(.A(G238), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n415), .A2(new_n418), .A3(new_n419), .A4(new_n320), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n410), .A2(new_n411), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n415), .A2(new_n418), .A3(new_n320), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT68), .A3(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(G200), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT12), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n264), .B2(new_n220), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n254), .A2(new_n220), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n268), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n359), .B2(new_n349), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n430), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT11), .B1(new_n430), .B2(new_n252), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n410), .A2(G190), .A3(new_n420), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n424), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n410), .A2(G179), .A3(new_n420), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n421), .A2(G169), .A3(new_n423), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n421), .A2(KEYINPUT14), .A3(G169), .A4(new_n423), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n435), .B1(new_n442), .B2(new_n433), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT69), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT69), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(new_n435), .C1(new_n442), .C2(new_n433), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n347), .B(new_n403), .C1(new_n444), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT81), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT80), .B1(new_n207), .B2(G107), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT23), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT23), .ZN(new_n451));
  OAI211_X1 g0251(.A(KEYINPUT80), .B(new_n451), .C1(new_n207), .C2(G107), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n450), .A2(new_n452), .B1(G116), .B2(new_n350), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  AOI21_X1  g0254(.A(G20), .B1(new_n276), .B2(new_n277), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G87), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n207), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT24), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(KEYINPUT22), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n296), .A2(new_n454), .A3(new_n207), .A4(G87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n453), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n348), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT73), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n206), .A2(G33), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n348), .A2(new_n467), .A3(new_n263), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n263), .A2(new_n468), .A3(new_n216), .A4(new_n251), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n471), .A3(G107), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n263), .A2(G107), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n448), .B1(new_n466), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n465), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n464), .B1(new_n463), .B2(new_n453), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n252), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n475), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT81), .ZN(new_n481));
  OAI211_X1 g0281(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n482));
  OAI211_X1 g0282(.A(G250), .B(new_n308), .C1(new_n270), .C2(new_n271), .ZN(new_n483));
  INV_X1    g0283(.A(G294), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n482), .B(new_n483), .C1(new_n275), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n306), .ZN(new_n486));
  INV_X1    g0286(.A(G45), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(G1), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT75), .ZN(new_n489));
  INV_X1    g0289(.A(G41), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(KEYINPUT75), .B2(G41), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n317), .A2(new_n488), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n488), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G264), .A3(new_n321), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n486), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G169), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n486), .A2(G179), .A3(new_n494), .A4(new_n496), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n476), .A2(new_n481), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n497), .A2(new_n337), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n497), .A2(G200), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n479), .A3(new_n480), .A4(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n505));
  OAI211_X1 g0305(.A(G257), .B(new_n308), .C1(new_n270), .C2(new_n271), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n306), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n495), .A2(G270), .A3(new_n321), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n494), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n470), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n264), .A2(new_n512), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n251), .A2(new_n216), .B1(G20), .B2(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n207), .C1(G33), .C2(new_n245), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT20), .B1(new_n515), .B2(new_n517), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n513), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n511), .A2(new_n520), .A3(G169), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n508), .A2(new_n306), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n510), .A2(new_n494), .ZN(new_n525));
  OAI21_X1  g0325(.A(G200), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n520), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n509), .A2(G190), .A3(new_n494), .A4(new_n510), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n524), .A2(new_n525), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G179), .A3(new_n520), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n511), .A2(new_n520), .A3(KEYINPUT21), .A4(G169), .ZN(new_n532));
  AND4_X1   g0332(.A1(new_n523), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n501), .A2(new_n504), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n207), .B(G68), .C1(new_n270), .C2(new_n271), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n349), .A2(new_n245), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(KEYINPUT19), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT77), .B(G87), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n538), .A2(new_n539), .B1(new_n207), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n252), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n385), .A2(new_n264), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n469), .A2(new_n471), .A3(G87), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n546));
  OAI211_X1 g0346(.A(G238), .B(new_n308), .C1(new_n270), .C2(new_n271), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n306), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n488), .A2(new_n223), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n321), .A2(new_n551), .B1(new_n317), .B2(new_n488), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(G190), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT78), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n206), .A2(G45), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n321), .A2(G250), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n321), .A2(G274), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(new_n555), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n306), .B2(new_n549), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n553), .B(new_n554), .C1(new_n340), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(KEYINPUT78), .A3(G190), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n545), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(G169), .B1(new_n550), .B2(new_n552), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n385), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n469), .A2(new_n471), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n542), .A2(new_n543), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n550), .A2(new_n323), .A3(new_n552), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT79), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT79), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n572));
  AND4_X1   g0372(.A1(KEYINPUT78), .A2(new_n550), .A3(G190), .A4(new_n552), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT78), .B1(new_n559), .B2(G190), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n550), .A2(new_n552), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n573), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n572), .C1(new_n577), .C2(new_n545), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(new_n308), .C1(new_n270), .C2(new_n271), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n296), .A2(KEYINPUT4), .A3(G244), .A4(new_n308), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n296), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n516), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n495), .A2(G257), .A3(new_n321), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n494), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT76), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n585), .A2(new_n306), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n494), .A3(KEYINPUT76), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n323), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n306), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n588), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n326), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n244), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g0397(.A(G97), .B(G107), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n268), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n207), .B1(new_n359), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n287), .A2(G107), .A3(new_n288), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT72), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n287), .A2(new_n288), .A3(KEYINPUT72), .A4(G107), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n348), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n608));
  OAI21_X1  g0408(.A(G97), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n264), .A2(G97), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(KEYINPUT74), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT74), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n245), .B1(new_n469), .B2(new_n471), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n610), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n591), .B(new_n595), .C1(new_n606), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n602), .A2(new_n603), .ZN(new_n618));
  INV_X1    g0418(.A(new_n601), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n605), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n252), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n612), .A2(new_n615), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n594), .A2(G200), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n589), .A2(G190), .A3(new_n590), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n534), .A2(new_n579), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n447), .A2(new_n627), .ZN(G372));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n291), .A2(new_n334), .A3(new_n331), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n334), .B1(new_n291), .B2(new_n331), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n333), .A2(KEYINPUT87), .A3(new_n335), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n343), .A2(new_n346), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n401), .A2(new_n400), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n435), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n442), .B2(new_n433), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n378), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n380), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n444), .A2(new_n446), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n403), .A2(new_n347), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT83), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT82), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n568), .B1(new_n563), .B2(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n559), .A2(KEYINPUT82), .A3(G169), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n563), .A2(new_n648), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT82), .B1(new_n559), .B2(G169), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT83), .A4(new_n568), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n567), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n621), .A2(new_n622), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT85), .ZN(new_n658));
  AOI21_X1  g0458(.A(G169), .B1(new_n589), .B2(new_n590), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n323), .A2(new_n592), .A3(new_n590), .A4(new_n593), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n620), .A2(new_n252), .B1(new_n615), .B2(new_n612), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n595), .A2(new_n591), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT85), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n577), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT84), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n545), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n545), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n656), .A2(new_n662), .A3(new_n665), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n663), .A2(new_n664), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n673), .A2(new_n570), .A3(new_n578), .ZN(new_n674));
  XNOR2_X1  g0474(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n646), .A2(new_n672), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n500), .B1(new_n466), .B2(new_n475), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n531), .A2(new_n532), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n523), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(new_n617), .A3(new_n625), .A4(new_n504), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n577), .B1(new_n669), .B2(new_n668), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n656), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n642), .B1(new_n645), .B2(new_n684), .ZN(G369));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n523), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n527), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n533), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n693), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n501), .A2(new_n692), .ZN(new_n699));
  INV_X1    g0499(.A(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n476), .A2(new_n481), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n501), .A2(new_n701), .A3(new_n504), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n501), .A2(new_n686), .A3(new_n504), .A4(new_n692), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n678), .A2(new_n700), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(G399));
  NAND2_X1  g0508(.A1(new_n210), .A2(new_n490), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n538), .A2(new_n512), .A3(new_n539), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n214), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT90), .B1(new_n672), .B2(new_n646), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n662), .A2(new_n665), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n682), .B1(new_n655), .B2(new_n567), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT26), .A4(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n675), .B1(new_n579), .B2(new_n617), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n715), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n617), .A2(new_n625), .A3(new_n504), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n523), .A2(new_n531), .A3(new_n532), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n501), .B2(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n724), .A2(new_n671), .B1(new_n567), .B2(new_n655), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n692), .B1(new_n677), .B2(new_n683), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n509), .A2(G179), .A3(new_n494), .A4(new_n510), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n486), .A2(new_n496), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n731), .A2(new_n732), .A3(new_n575), .ZN(new_n733));
  INV_X1    g0533(.A(new_n594), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(KEYINPUT89), .A2(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n530), .A2(G179), .A3(new_n559), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n594), .A3(new_n497), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n733), .B(new_n734), .C1(KEYINPUT89), .C2(KEYINPUT30), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n627), .B2(new_n692), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n700), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n742), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n727), .A2(new_n730), .B1(G330), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n714), .B1(new_n748), .B2(G1), .ZN(G364));
  INV_X1    g0549(.A(new_n709), .ZN(new_n750));
  INV_X1    g0550(.A(G13), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n206), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n210), .A2(new_n296), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n210), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n242), .A2(new_n487), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n210), .A2(new_n272), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n487), .B2(new_n215), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n216), .B1(G20), .B2(new_n326), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n755), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n323), .A2(new_n340), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G294), .ZN(new_n774));
  NAND3_X1  g0574(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(G317), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT33), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT33), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n207), .A2(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n323), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n780), .B(new_n272), .C1(new_n781), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n775), .A2(new_n337), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(G326), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n771), .A2(new_n782), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G303), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(new_n337), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n340), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n783), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n791), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n782), .A2(new_n793), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(G283), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n774), .A2(new_n787), .A3(new_n790), .A4(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n795), .A2(new_n266), .B1(new_n784), .B2(new_n359), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G50), .B2(new_n786), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT92), .Z(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n788), .A2(KEYINPUT32), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n773), .A2(G97), .ZN(new_n807));
  INV_X1    g0607(.A(new_n776), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n220), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n794), .A2(new_n538), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n798), .A2(new_n243), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n272), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n788), .B2(new_n805), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n806), .A2(new_n807), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n801), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n769), .B1(new_n815), .B2(new_n766), .ZN(new_n816));
  INV_X1    g0616(.A(new_n765), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n696), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT91), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n697), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n696), .A2(KEYINPUT91), .A3(G330), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n755), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n696), .B2(G330), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n818), .B1(new_n822), .B2(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n395), .A2(new_n399), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n700), .A2(new_n388), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n636), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n636), .A2(new_n692), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n692), .B(new_n831), .C1(new_n677), .C2(new_n683), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n672), .A2(new_n646), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n674), .A2(new_n676), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n683), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n700), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT96), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n826), .A2(new_n827), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n838), .B(new_n829), .C1(new_n839), .C2(new_n636), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT96), .B1(new_n828), .B2(new_n830), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n832), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n747), .A2(G330), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n755), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n766), .A2(new_n763), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n755), .B1(G77), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n272), .B1(new_n794), .B2(new_n243), .C1(new_n851), .C2(new_n808), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G303), .B2(new_n786), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n789), .A2(G311), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n795), .A2(new_n484), .B1(new_n784), .B2(new_n512), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G87), .B2(new_n799), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n853), .A2(new_n807), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n795), .ZN(new_n858));
  INV_X1    g0658(.A(new_n784), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G143), .A2(new_n858), .B1(new_n859), .B2(G159), .ZN(new_n860));
  INV_X1    g0660(.A(new_n786), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  INV_X1    g0662(.A(G150), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n860), .B1(new_n861), .B2(new_n862), .C1(new_n863), .C2(new_n808), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n773), .A2(new_n260), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n296), .B1(new_n798), .B2(new_n220), .C1(new_n202), .C2(new_n794), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n789), .B2(G132), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n864), .A2(new_n865), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n857), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n850), .B1(new_n872), .B2(new_n766), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT94), .Z(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n764), .B2(new_n831), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT95), .Z(new_n876));
  NOR2_X1   g0676(.A1(new_n847), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(G384));
  NOR2_X1   g0678(.A1(new_n752), .A2(new_n206), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n690), .B(KEYINPUT88), .Z(new_n881));
  INV_X1    g0681(.A(KEYINPUT16), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n201), .B1(new_n260), .B2(G68), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n883), .A2(new_n207), .B1(new_n805), .B2(new_n600), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n220), .B1(new_n285), .B2(new_n278), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n281), .A3(new_n252), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n881), .B1(new_n887), .B2(new_n265), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n347), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n291), .A2(new_n691), .ZN(new_n890));
  XNOR2_X1  g0690(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n332), .A2(new_n890), .A3(new_n344), .A4(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n344), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n265), .A2(new_n887), .B1(new_n330), .B2(new_n881), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT100), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(KEYINPUT38), .B(new_n889), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n742), .A2(KEYINPUT102), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n741), .A2(new_n905), .A3(KEYINPUT31), .A4(new_n700), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n744), .B2(new_n746), .ZN(new_n909));
  INV_X1    g0709(.A(new_n831), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n440), .A2(new_n441), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n436), .ZN(new_n912));
  INV_X1    g0712(.A(new_n433), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT97), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT97), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n442), .B2(new_n433), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n692), .A2(new_n433), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n917), .A2(KEYINPUT98), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(KEYINPUT98), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n918), .A2(new_n435), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n914), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n442), .A2(new_n435), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n917), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n910), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n903), .A2(new_n909), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n926));
  INV_X1    g0726(.A(new_n890), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n332), .A2(new_n890), .A3(new_n344), .ZN(new_n929));
  INV_X1    g0729(.A(new_n891), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n892), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n900), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n880), .B1(new_n934), .B2(new_n902), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n921), .A2(new_n923), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n831), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n501), .A2(new_n504), .A3(new_n533), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n570), .A2(new_n578), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n617), .A2(new_n625), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n692), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT31), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n907), .B1(new_n942), .B2(new_n745), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n880), .A2(new_n925), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n946), .A2(new_n645), .A3(new_n943), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n447), .B2(new_n909), .ZN(new_n948));
  INV_X1    g0748(.A(G330), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT103), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n729), .B(new_n700), .C1(new_n721), .C2(new_n725), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n447), .B1(new_n837), .B2(KEYINPUT29), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT101), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n645), .B1(new_n729), .B2(new_n728), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT101), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n727), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n641), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n926), .A2(new_n927), .B1(new_n892), .B2(new_n931), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n902), .B1(new_n959), .B2(KEYINPUT38), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT39), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n914), .A2(new_n916), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n700), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n902), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n832), .A2(new_n829), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n903), .A3(new_n936), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n634), .A2(new_n881), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n958), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n879), .B1(new_n951), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n951), .B2(new_n972), .ZN(new_n974));
  INV_X1    g0774(.A(new_n599), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT35), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT35), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(G116), .A3(new_n217), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT36), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n215), .B(G77), .C1(new_n220), .C2(new_n266), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(G50), .B2(new_n220), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(G1), .A3(new_n751), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n974), .A2(new_n979), .A3(new_n982), .ZN(G367));
  OAI211_X1 g0783(.A(new_n617), .B(new_n625), .C1(new_n663), .C2(new_n692), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n617), .B1(new_n984), .B2(new_n501), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n692), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n673), .A2(new_n700), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(new_n705), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT42), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n700), .A2(new_n669), .A3(new_n668), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n656), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n718), .B2(new_n994), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  AOI211_X1 g0798(.A(KEYINPUT43), .B(new_n995), .C1(new_n718), .C2(new_n994), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n986), .C1(new_n991), .C2(new_n992), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT104), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(KEYINPUT104), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n704), .A2(new_n988), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n705), .A2(new_n706), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT105), .B1(new_n988), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT105), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n984), .A2(new_n987), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n707), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT44), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n707), .B2(new_n1010), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n988), .A2(KEYINPUT44), .A3(new_n1007), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1012), .A2(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1008), .A2(new_n1011), .A3(KEYINPUT45), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n1017), .A2(new_n704), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n704), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n699), .B(new_n702), .C1(new_n723), .C2(new_n700), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n705), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n820), .A3(new_n821), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n698), .A2(new_n705), .A3(new_n1022), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n837), .A2(KEYINPUT29), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n844), .C1(new_n952), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1021), .A2(KEYINPUT106), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT106), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1018), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n704), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1017), .A2(new_n704), .A3(new_n1018), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1032), .B1(new_n1039), .B2(new_n1029), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1031), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1006), .B1(new_n1041), .B2(new_n748), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1005), .B1(new_n1042), .B2(new_n754), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G97), .A2(new_n799), .B1(new_n859), .B2(G283), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n296), .B1(new_n858), .B2(G303), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n777), .C2(new_n788), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n794), .A2(new_n512), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT46), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n484), .B2(new_n808), .C1(new_n781), .C2(new_n861), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1046), .B(new_n1050), .C1(G107), .C2(new_n773), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n773), .A2(G68), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n858), .A2(G150), .B1(G143), .B2(new_n786), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT107), .Z(new_n1055));
  INV_X1    g0855(.A(new_n794), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1056), .A2(new_n260), .B1(new_n859), .B2(G50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n272), .B1(new_n799), .B2(G77), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n805), .C2(new_n808), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G137), .B2(new_n789), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1051), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n766), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n767), .B1(new_n210), .B2(new_n385), .C1(new_n238), .C2(new_n760), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n755), .A3(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n996), .A2(new_n765), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1043), .A2(new_n1069), .ZN(G387));
  NOR2_X1   g0870(.A1(new_n861), .A2(new_n805), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n272), .B1(new_n799), .B2(G97), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n202), .B2(new_n795), .C1(new_n359), .C2(new_n794), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT110), .B(G150), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1071), .B(new_n1073), .C1(new_n789), .C2(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n261), .A2(new_n776), .B1(new_n859), .B2(G68), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT111), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n773), .A2(new_n565), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n789), .A2(G326), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n296), .B1(new_n799), .B2(G116), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n795), .A2(new_n777), .B1(new_n784), .B2(new_n791), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT112), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n808), .A2(new_n781), .B1(new_n861), .B2(new_n796), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT48), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(KEYINPUT48), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n773), .A2(G283), .B1(G294), .B2(new_n1056), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT113), .Z(new_n1092));
  INV_X1    g0892(.A(KEYINPUT49), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1080), .B(new_n1081), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1079), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n766), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n235), .A2(G45), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT109), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n383), .A2(new_n202), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT50), .Z(new_n1101));
  AOI211_X1 g0901(.A(G45), .B(new_n710), .C1(G68), .C2(G77), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n760), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(G107), .B2(new_n210), .C1(new_n711), .C2(new_n756), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n823), .B1(new_n1105), .B2(new_n767), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1097), .B(new_n1106), .C1(new_n703), .C2(new_n817), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1029), .A2(new_n750), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n748), .A2(new_n1027), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1107), .B1(new_n753), .B2(new_n1026), .C1(new_n1108), .C2(new_n1109), .ZN(G393));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1037), .A2(new_n1111), .A3(new_n1038), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1035), .A2(KEYINPUT114), .A3(new_n1036), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n988), .A2(new_n765), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n767), .B1(new_n245), .B2(new_n210), .C1(new_n249), .C2(new_n760), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n755), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n296), .B1(new_n798), .B2(new_n222), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n383), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1119), .A2(new_n784), .B1(new_n220), .B2(new_n794), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(G50), .C2(new_n776), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n861), .A2(new_n863), .B1(new_n795), .B2(new_n805), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n773), .A2(G77), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n789), .A2(G143), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n859), .A2(G294), .B1(G303), .B2(new_n776), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n773), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n512), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT116), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n861), .A2(new_n777), .B1(new_n795), .B2(new_n781), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT52), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n296), .B(new_n811), .C1(G283), .C2(new_n1056), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n796), .C2(new_n788), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1127), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1117), .B1(new_n1136), .B2(new_n766), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1114), .A2(new_n754), .B1(new_n1115), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1041), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n750), .B1(new_n1114), .B2(new_n1030), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(G390));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n909), .A2(new_n924), .A3(G330), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n964), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n960), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n700), .B1(new_n721), .B2(new_n725), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n828), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n829), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1146), .B1(new_n1150), .B2(new_n936), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n967), .A2(new_n936), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1152), .A2(new_n1145), .B1(new_n962), .B2(new_n965), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1144), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1145), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n962), .A2(new_n965), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n830), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n936), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n960), .B(new_n1145), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n747), .A2(G330), .A3(new_n831), .A4(new_n936), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1157), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1156), .A2(new_n763), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n858), .A2(G132), .B1(new_n859), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n272), .B1(new_n799), .B2(G50), .ZN(new_n1168));
  INV_X1    g0968(.A(G125), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1168), .C1(new_n1169), .C2(new_n788), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1056), .A2(new_n1074), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n861), .C1(new_n862), .C2(new_n808), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1170), .B(new_n1175), .C1(G159), .C2(new_n773), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n296), .B1(new_n799), .B2(G68), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n861), .B2(new_n851), .C1(new_n243), .C2(new_n808), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G87), .A2(new_n1056), .B1(new_n858), .B2(G116), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n245), .B2(new_n784), .C1(new_n484), .C2(new_n788), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G77), .C2(new_n773), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n766), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n755), .C1(new_n261), .C2(new_n849), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT119), .Z(new_n1184));
  AOI22_X1  g0984(.A1(new_n1163), .A2(new_n754), .B1(new_n1164), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT117), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n967), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n746), .B1(new_n941), .B2(KEYINPUT31), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n742), .ZN(new_n1189));
  OAI211_X1 g0989(.A(G330), .B(new_n831), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1159), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1187), .B1(new_n1191), .B2(new_n1143), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n842), .B(G330), .C1(new_n1188), .C2(new_n907), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1159), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1192), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n909), .A2(G330), .A3(new_n447), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n955), .A2(new_n727), .A3(new_n956), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n956), .B1(new_n955), .B2(new_n727), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n642), .B(new_n1197), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1186), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1158), .A2(new_n1161), .A3(new_n1195), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n944), .A2(G330), .B1(new_n1159), .B2(new_n1190), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n1187), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1205), .A2(new_n958), .A3(KEYINPUT117), .A4(new_n1197), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n750), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1202), .B1(new_n1201), .B2(new_n1206), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1142), .B(new_n1185), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1197), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n641), .B(new_n1212), .C1(new_n954), .C2(new_n957), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT117), .B1(new_n1213), .B2(new_n1205), .ZN(new_n1214));
  AND4_X1   g1014(.A1(KEYINPUT117), .A2(new_n1205), .A3(new_n958), .A4(new_n1197), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1163), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n750), .A3(new_n1207), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1142), .B1(new_n1217), .B2(new_n1185), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1211), .A2(new_n1218), .ZN(G378));
  NAND2_X1  g1019(.A1(new_n378), .A2(new_n380), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n691), .B1(new_n353), .B2(new_n355), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1220), .B(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n763), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n755), .B1(G50), .B2(new_n849), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n275), .A2(new_n490), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT121), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n202), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n490), .B2(new_n272), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G41), .B(new_n296), .C1(new_n1056), .C2(G77), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n245), .B2(new_n808), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G116), .B2(new_n786), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n799), .A2(new_n260), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n243), .B2(new_n795), .C1(new_n385), .C2(new_n784), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G283), .B2(new_n789), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1237), .A3(new_n1052), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT58), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1174), .A2(new_n795), .B1(new_n794), .B2(new_n1165), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G137), .B2(new_n859), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G125), .A2(new_n786), .B1(new_n776), .B2(G132), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(new_n1129), .C2(new_n863), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n798), .A2(new_n805), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1229), .B(new_n1247), .C1(new_n789), .C2(G124), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1240), .B1(new_n1239), .B2(new_n1238), .C1(new_n1245), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1227), .B1(new_n1250), .B2(new_n766), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1224), .B1(new_n945), .B2(G330), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n936), .B(new_n831), .C1(new_n1188), .C2(new_n907), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n892), .A2(new_n895), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT100), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT38), .B1(new_n1259), .B2(new_n889), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n902), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n880), .B1(new_n1255), .B2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n909), .A2(new_n960), .A3(new_n924), .A4(KEYINPUT40), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(G330), .A3(new_n1264), .A4(new_n1224), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n970), .B1(new_n1254), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(G330), .A3(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1225), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n971), .A3(new_n1265), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT122), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1267), .A2(KEYINPUT122), .A3(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1253), .B1(new_n1275), .B2(new_n754), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1216), .A2(new_n1213), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1275), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1200), .B1(new_n1279), .B2(new_n1163), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1271), .A2(KEYINPUT57), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n750), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1276), .B1(new_n1278), .B2(new_n1282), .ZN(G375));
  NAND2_X1  g1083(.A1(new_n1159), .A2(new_n763), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n755), .B1(G68), .B2(new_n849), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G137), .A2(new_n858), .B1(new_n859), .B2(G150), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n805), .B2(new_n794), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G128), .B2(new_n789), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1235), .B(new_n296), .C1(new_n808), .C2(new_n1165), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(G132), .B2(new_n786), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1288), .B(new_n1290), .C1(new_n202), .C2(new_n1129), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n272), .B1(new_n798), .B2(new_n359), .C1(new_n861), .C2(new_n484), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(G116), .B2(new_n776), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n789), .A2(G303), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n795), .A2(new_n851), .B1(new_n784), .B2(new_n243), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G97), .B2(new_n1056), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1078), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1285), .B1(new_n1298), .B2(new_n766), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1205), .A2(new_n754), .B1(new_n1284), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT123), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1196), .A2(new_n1200), .A3(KEYINPUT123), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1006), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1201), .A2(new_n1306), .A3(new_n1206), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1305), .B2(new_n1307), .ZN(G381));
  OAI21_X1  g1108(.A(new_n1185), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1309));
  OR2_X1    g1109(.A1(G393), .A2(G396), .ZN(new_n1310));
  OR4_X1    g1110(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1310), .ZN(new_n1311));
  OR4_X1    g1111(.A1(new_n1309), .A2(new_n1311), .A3(G375), .A4(G381), .ZN(G407));
  AND3_X1   g1112(.A1(new_n1269), .A2(new_n971), .A3(new_n1265), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n971), .B1(new_n1269), .B2(new_n1265), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1272), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT122), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n754), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1252), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1281), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n709), .B1(new_n1277), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT57), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1321), .B1(new_n1322), .B2(new_n1280), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1318), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1309), .ZN(new_n1325));
  INV_X1    g1125(.A(G343), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(G213), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(KEYINPUT124), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1324), .A2(new_n1325), .A3(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(G407), .A2(G213), .A3(new_n1329), .ZN(G409));
  INV_X1    g1130(.A(KEYINPUT60), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n750), .B1(new_n1301), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1201), .A2(KEYINPUT60), .A3(new_n1206), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1333), .B1(new_n1334), .B2(new_n1305), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(G384), .A3(new_n1300), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1196), .A2(new_n1200), .A3(KEYINPUT123), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT123), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1201), .A2(KEYINPUT60), .A3(new_n1206), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1332), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1300), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n877), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1327), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(G2897), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1336), .A2(new_n1343), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1328), .A2(G2897), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1347), .B1(new_n1336), .B2(new_n1343), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1277), .A2(new_n1275), .A3(new_n1306), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1253), .B1(new_n1271), .B2(new_n754), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1309), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1352), .B1(G378), .B2(new_n1324), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1349), .B1(new_n1353), .B2(new_n1344), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1325), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1309), .A2(KEYINPUT120), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n1210), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1356), .B1(G375), .B2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1328), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1336), .A2(new_n1343), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT63), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1359), .A2(new_n1360), .A3(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT106), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1039), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n748), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n754), .B1(new_n1367), .B2(new_n1306), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1004), .ZN(new_n1369));
  XNOR2_X1  g1169(.A(new_n1003), .B(new_n1369), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1069), .B(G390), .C1(new_n1368), .C2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(KEYINPUT126), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT125), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(G390), .A2(new_n1373), .ZN(new_n1374));
  OAI211_X1 g1174(.A(KEYINPUT125), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1367), .A2(new_n1306), .ZN(new_n1376));
  AOI21_X1  g1176(.A(new_n1370), .B1(new_n1376), .B2(new_n753), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1374), .B(new_n1375), .C1(new_n1377), .C2(new_n1068), .ZN(new_n1378));
  XOR2_X1   g1178(.A(G393), .B(G396), .Z(new_n1379));
  INV_X1    g1179(.A(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT126), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1043), .A2(new_n1381), .A3(new_n1069), .A4(G390), .ZN(new_n1382));
  NAND4_X1  g1182(.A1(new_n1372), .A2(new_n1378), .A3(new_n1380), .A4(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1371), .ZN(new_n1384));
  AOI21_X1  g1184(.A(G390), .B1(new_n1043), .B2(new_n1069), .ZN(new_n1385));
  OAI21_X1  g1185(.A(new_n1379), .B1(new_n1384), .B2(new_n1385), .ZN(new_n1386));
  AOI21_X1  g1186(.A(KEYINPUT61), .B1(new_n1383), .B2(new_n1386), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1354), .A2(new_n1364), .A3(new_n1387), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(G378), .A2(new_n1324), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1344), .B1(new_n1389), .B2(new_n1356), .ZN(new_n1390));
  INV_X1    g1190(.A(new_n1361), .ZN(new_n1391));
  AOI21_X1  g1191(.A(KEYINPUT63), .B1(new_n1390), .B2(new_n1391), .ZN(new_n1392));
  OAI21_X1  g1192(.A(KEYINPUT127), .B1(new_n1388), .B2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1383), .A2(new_n1386), .ZN(new_n1394));
  INV_X1    g1194(.A(KEYINPUT61), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1359), .A2(new_n1327), .ZN(new_n1397));
  AOI21_X1  g1197(.A(new_n1396), .B1(new_n1397), .B2(new_n1349), .ZN(new_n1398));
  INV_X1    g1198(.A(KEYINPUT127), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1359), .A2(new_n1327), .A3(new_n1391), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1400), .A2(new_n1362), .ZN(new_n1401));
  NAND4_X1  g1201(.A1(new_n1398), .A2(new_n1399), .A3(new_n1401), .A4(new_n1364), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1393), .A2(new_n1402), .ZN(new_n1403));
  INV_X1    g1203(.A(new_n1394), .ZN(new_n1404));
  INV_X1    g1204(.A(KEYINPUT62), .ZN(new_n1405));
  NOR2_X1   g1205(.A1(new_n1353), .A2(new_n1328), .ZN(new_n1406));
  NOR2_X1   g1206(.A1(new_n1361), .A2(new_n1405), .ZN(new_n1407));
  AOI22_X1  g1207(.A1(new_n1405), .A2(new_n1400), .B1(new_n1406), .B2(new_n1407), .ZN(new_n1408));
  OAI21_X1  g1208(.A(new_n1349), .B1(new_n1353), .B2(new_n1328), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1409), .A2(new_n1395), .ZN(new_n1410));
  OAI21_X1  g1210(.A(new_n1404), .B1(new_n1408), .B2(new_n1410), .ZN(new_n1411));
  NAND2_X1  g1211(.A1(new_n1403), .A2(new_n1411), .ZN(G405));
  NAND2_X1  g1212(.A1(G375), .A2(new_n1325), .ZN(new_n1413));
  AND2_X1   g1213(.A1(new_n1389), .A2(new_n1413), .ZN(new_n1414));
  OR2_X1    g1214(.A1(new_n1414), .A2(new_n1361), .ZN(new_n1415));
  NAND2_X1  g1215(.A1(new_n1414), .A2(new_n1361), .ZN(new_n1416));
  AND3_X1   g1216(.A1(new_n1415), .A2(new_n1416), .A3(new_n1404), .ZN(new_n1417));
  AOI21_X1  g1217(.A(new_n1404), .B1(new_n1415), .B2(new_n1416), .ZN(new_n1418));
  NOR2_X1   g1218(.A1(new_n1417), .A2(new_n1418), .ZN(G402));
endmodule


