//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G238), .Z(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n202), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n217), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n209), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT7), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT7), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n252), .A2(new_n256), .A3(new_n209), .A4(new_n253), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G68), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT16), .ZN(new_n259));
  XNOR2_X1  g0059(.A(G58), .B(G68), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n260), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n258), .B2(new_n262), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n249), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n249), .B1(new_n208), .B2(G20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(new_n267), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT70), .B1(new_n265), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT18), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G232), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(G223), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n288), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G87), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n282), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n298), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  INV_X1    g0103(.A(new_n249), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n258), .A2(new_n262), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT16), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n271), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n271), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(new_n301), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT71), .A2(KEYINPUT18), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n275), .A2(new_n276), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n287), .B2(new_n297), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n282), .B1(new_n293), .B2(new_n294), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n319), .A2(KEYINPUT72), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(KEYINPUT72), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n318), .A2(new_n286), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT17), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n265), .A2(new_n324), .A3(new_n271), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n302), .A2(new_n315), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n331));
  INV_X1    g0131(.A(G150), .ZN(new_n332));
  INV_X1    g0132(.A(new_n261), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n209), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n266), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n249), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n270), .A2(G50), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(G50), .C2(new_n268), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT9), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n280), .B1(new_n284), .B2(new_n289), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n291), .A2(new_n292), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT65), .B(G223), .Z(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G1698), .ZN(new_n345));
  OR2_X1    g0145(.A1(G222), .A2(G1698), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n252), .A2(new_n253), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n296), .B1(new_n348), .B2(G77), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n319), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT66), .B(G200), .Z(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(new_n350), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n340), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT10), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(KEYINPUT10), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n280), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n282), .A2(G244), .A3(new_n283), .ZN(new_n361));
  INV_X1    g0161(.A(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n348), .A2(G232), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G107), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n348), .A2(G1698), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n363), .B1(new_n364), .B2(new_n348), .C1(new_n365), .C2(new_n220), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n360), .B(new_n361), .C1(new_n366), .C2(new_n296), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n367), .A2(new_n300), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n270), .A2(G77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G20), .A2(G77), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n335), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n261), .B2(new_n267), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n369), .B1(G77), .B2(new_n268), .C1(new_n373), .C2(new_n304), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n367), .B2(G169), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n367), .B2(G190), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n352), .B2(new_n367), .ZN(new_n379));
  INV_X1    g0179(.A(new_n350), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n339), .B1(new_n380), .B2(G169), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n350), .A2(G179), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  OR3_X1    g0184(.A1(new_n330), .A2(new_n359), .A3(new_n384), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n333), .A2(new_n241), .B1(new_n209), .B2(G68), .ZN(new_n386));
  INV_X1    g0186(.A(G77), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n335), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n249), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n270), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT12), .ZN(new_n393));
  INV_X1    g0193(.A(new_n268), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n202), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n392), .A2(new_n202), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n389), .A2(new_n390), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n391), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n282), .A2(G238), .A3(new_n283), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n280), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT68), .ZN(new_n404));
  OAI211_X1 g0204(.A(G226), .B(new_n362), .C1(new_n291), .C2(new_n292), .ZN(new_n405));
  OAI211_X1 g0205(.A(G232), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G97), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT67), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT67), .A4(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n296), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n404), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n401), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n416), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n417), .A2(new_n418), .B1(new_n419), .B2(new_n300), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n418), .A3(G169), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n400), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT69), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(new_n399), .C1(new_n319), .C2(new_n419), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n423), .B2(new_n426), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n385), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT5), .B(G41), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n208), .A2(G45), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n217), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n430), .A2(new_n432), .B1(new_n433), .B2(new_n281), .ZN(new_n434));
  OR2_X1    g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G274), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n433), .B2(new_n281), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n434), .A2(G270), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n441));
  OAI211_X1 g0241(.A(G257), .B(new_n362), .C1(new_n291), .C2(new_n292), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n252), .A2(G303), .A3(new_n253), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n296), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n445), .A3(G179), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n268), .A2(G116), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n208), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n268), .A2(new_n449), .A3(new_n217), .A4(new_n248), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT20), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n209), .B1(new_n454), .B2(G33), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT75), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT75), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G33), .A3(G283), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n248), .A2(new_n217), .B1(G20), .B2(new_n451), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n453), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n457), .A2(new_n459), .ZN(new_n464));
  OAI211_X1 g0264(.A(KEYINPUT20), .B(new_n461), .C1(new_n464), .C2(new_n455), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n452), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n446), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n465), .ZN(new_n468));
  INV_X1    g0268(.A(new_n452), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n401), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n444), .A2(new_n296), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n430), .A2(new_n432), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G270), .A3(new_n282), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n437), .A2(new_n439), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT80), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT80), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n440), .A2(new_n445), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n467), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n440), .A2(new_n477), .A3(new_n445), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n477), .B1(new_n440), .B2(new_n445), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n482), .A2(new_n483), .B1(new_n320), .B2(new_n321), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n476), .A2(G200), .A3(new_n478), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(new_n466), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n482), .A2(new_n483), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT21), .A3(new_n470), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n481), .A2(new_n486), .A3(new_n488), .A4(KEYINPUT81), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(G244), .B(new_n362), .C1(new_n291), .C2(new_n292), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n348), .A2(KEYINPUT4), .A3(G244), .A4(new_n362), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n457), .A2(new_n459), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n348), .A2(G250), .A3(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n500), .A2(new_n296), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n434), .A2(G257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n474), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n401), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n500), .A2(new_n506), .A3(new_n296), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n500), .B2(new_n296), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n300), .B(new_n505), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT77), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT74), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT6), .ZN(new_n512));
  AND2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n205), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n364), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n209), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n333), .A2(new_n387), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n517), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n364), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  XNOR2_X1  g0320(.A(G97), .B(G107), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(new_n512), .ZN(new_n522));
  OAI211_X1 g0322(.A(KEYINPUT74), .B(new_n519), .C1(new_n522), .C2(new_n209), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n255), .A2(G107), .A3(new_n257), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n249), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n394), .A2(new_n454), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n450), .B2(new_n454), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n510), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AOI211_X1 g0330(.A(KEYINPUT77), .B(new_n528), .C1(new_n525), .C2(new_n249), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n504), .B(new_n509), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n528), .B1(new_n525), .B2(new_n249), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n503), .B1(new_n296), .B2(new_n500), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n431), .A2(G250), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n296), .A2(new_n539), .B1(new_n438), .B2(new_n431), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G238), .B(new_n362), .C1(new_n291), .C2(new_n292), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n348), .A2(KEYINPUT78), .A3(G244), .A4(G1698), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n296), .B1(new_n549), .B2(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  INV_X1    g0351(.A(new_n544), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n551), .A2(KEYINPUT79), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n300), .B(new_n541), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n371), .A2(new_n394), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n348), .A2(new_n209), .A3(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n209), .B1(new_n407), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G87), .B2(new_n206), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n335), .B2(new_n454), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n555), .B1(new_n561), .B2(new_n304), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n450), .A2(new_n371), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n551), .A2(new_n552), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n282), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n549), .A2(KEYINPUT79), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n540), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n554), .B(new_n565), .C1(new_n570), .C2(G169), .ZN(new_n571));
  INV_X1    g0371(.A(new_n450), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n562), .B1(G87), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G190), .B(new_n541), .C1(new_n550), .C2(new_n553), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n570), .C2(new_n352), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n532), .A2(new_n538), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n209), .A3(G87), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n343), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n543), .A2(G20), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT23), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n209), .B2(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n364), .A2(KEYINPUT23), .A3(G20), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G87), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(KEYINPUT82), .A3(G20), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n348), .A2(KEYINPUT22), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n580), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n580), .A2(new_n588), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n304), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n394), .A2(KEYINPUT25), .A3(new_n364), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT25), .B1(new_n394), .B2(new_n364), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(new_n364), .B2(new_n450), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n598));
  OAI211_X1 g0398(.A(G250), .B(new_n362), .C1(new_n291), .C2(new_n292), .ZN(new_n599));
  INV_X1    g0399(.A(G294), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n251), .C2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n296), .B1(G264), .B2(new_n434), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n474), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n597), .B(new_n604), .C1(new_n319), .C2(new_n603), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n401), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n300), .A3(new_n474), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n593), .C2(new_n596), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n429), .A2(new_n493), .A3(new_n576), .A4(new_n609), .ZN(new_n610));
  XOR2_X1   g0410(.A(new_n610), .B(KEYINPUT83), .Z(G372));
  INV_X1    g0411(.A(new_n383), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n265), .A2(new_n271), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n301), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT18), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n276), .A3(new_n301), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n423), .A2(new_n377), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n426), .A2(new_n329), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n357), .B2(new_n358), .ZN(new_n622));
  INV_X1    g0422(.A(new_n358), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(KEYINPUT85), .A3(new_n356), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n612), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n429), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n575), .A2(new_n571), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n628), .B2(new_n532), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n526), .A2(new_n529), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n509), .A2(new_n630), .A3(new_n504), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n571), .A3(new_n575), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(KEYINPUT26), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n541), .B1(new_n550), .B2(new_n553), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n564), .B1(new_n636), .B2(new_n401), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n635), .B1(new_n637), .B2(new_n554), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n532), .A2(new_n538), .A3(new_n571), .A4(new_n575), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n481), .A2(new_n488), .A3(new_n608), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n605), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n626), .B1(new_n627), .B2(new_n645), .ZN(G369));
  NAND2_X1  g0446(.A1(new_n481), .A2(new_n488), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n466), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n493), .A2(KEYINPUT86), .B1(new_n466), .B2(new_n654), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n493), .A2(KEYINPUT86), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n608), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n653), .B1(new_n593), .B2(new_n596), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n605), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n608), .A2(new_n653), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n647), .A2(new_n654), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n212), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n215), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n644), .A2(new_n654), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT90), .B1(new_n634), .B2(new_n638), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n509), .A2(new_n504), .ZN(new_n688));
  INV_X1    g0488(.A(new_n530), .ZN(new_n689));
  INV_X1    g0489(.A(new_n531), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n571), .A4(new_n575), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n687), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT90), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n637), .A2(new_n635), .A3(new_n554), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n640), .B2(new_n642), .ZN(new_n700));
  OAI211_X1 g0500(.A(KEYINPUT29), .B(new_n654), .C1(new_n695), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n686), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT89), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n446), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n704), .A2(new_n536), .A3(new_n602), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n440), .A2(new_n445), .A3(KEYINPUT89), .A4(G179), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n570), .A4(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n704), .A2(new_n536), .A3(new_n602), .A4(new_n706), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n636), .ZN(new_n710));
  AOI21_X1  g0510(.A(G179), .B1(new_n602), .B2(new_n474), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n533), .A2(new_n636), .A3(new_n487), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n713), .B2(new_n653), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n493), .A2(new_n576), .A3(new_n609), .A4(new_n654), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n702), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n683), .B1(new_n721), .B2(G1), .ZN(G364));
  NAND2_X1  g0522(.A1(new_n209), .A2(G13), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT91), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G45), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G1), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n678), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n660), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n659), .ZN(new_n729));
  INV_X1    g0529(.A(new_n727), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n677), .A2(new_n343), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n451), .B2(new_n677), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n677), .A2(new_n348), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G45), .B2(new_n215), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n246), .A2(new_n278), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n217), .B1(G20), .B2(new_n401), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n730), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  INV_X1    g0543(.A(new_n740), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n209), .A2(new_n300), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT33), .B(G317), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n750), .A2(KEYINPUT95), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(KEYINPUT95), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n748), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n209), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n353), .A2(new_n319), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(G283), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n353), .A2(G190), .A3(new_n754), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n322), .A2(new_n746), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G326), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n319), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n209), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n762), .A2(new_n763), .B1(new_n600), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(KEYINPUT94), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(KEYINPUT94), .ZN(new_n768));
  NOR4_X1   g0568(.A1(new_n209), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n348), .B1(new_n769), .B2(G329), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n745), .A2(new_n316), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n322), .A2(new_n771), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n770), .B1(new_n773), .B2(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OR4_X1    g0578(.A1(new_n760), .A2(new_n767), .A3(new_n768), .A4(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n201), .B1(new_n773), .B2(new_n387), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT93), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n348), .B1(new_n762), .B2(new_n241), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n755), .A2(new_n364), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n759), .A2(new_n586), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n780), .A2(new_n781), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n748), .A2(new_n202), .B1(new_n765), .B2(new_n454), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n769), .A2(G159), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n782), .A2(new_n786), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n739), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n743), .B1(new_n744), .B2(new_n793), .C1(new_n659), .C2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n729), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n374), .A2(new_n653), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n379), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n377), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n376), .A2(new_n654), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n684), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n802), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n654), .B(new_n805), .C1(new_n633), .C2(new_n643), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n727), .B1(new_n807), .B2(new_n719), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n719), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n740), .A2(new_n737), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT96), .Z(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n730), .B1(new_n387), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n756), .A2(G87), .ZN(new_n814));
  INV_X1    g0614(.A(new_n769), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n774), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(KEYINPUT98), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(KEYINPUT98), .ZN(new_n819));
  INV_X1    g0619(.A(new_n765), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n348), .B1(new_n820), .B2(G97), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n759), .B2(new_n364), .C1(new_n600), .C2(new_n776), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G116), .A2(new_n772), .B1(new_n747), .B2(G283), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n758), .B2(new_n762), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT97), .Z(new_n826));
  AOI22_X1  g0626(.A1(new_n761), .A2(G137), .B1(new_n747), .B2(G150), .ZN(new_n827));
  INV_X1    g0627(.A(G143), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(new_n828), .B2(new_n776), .C1(new_n829), .C2(new_n773), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n348), .B1(new_n815), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G58), .B2(new_n820), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n241), .B2(new_n759), .C1(new_n202), .C2(new_n755), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n831), .B2(KEYINPUT34), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n823), .A2(new_n826), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n813), .B1(new_n744), .B2(new_n838), .C1(new_n805), .C2(new_n738), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n809), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  INV_X1    g0641(.A(new_n522), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(KEYINPUT35), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(KEYINPUT35), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(G116), .A4(new_n218), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT36), .Z(new_n846));
  OAI211_X1 g0646(.A(new_n216), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n208), .B(G13), .C1(new_n847), .C2(new_n242), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n686), .A2(new_n429), .A3(new_n701), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n626), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT102), .ZN(new_n852));
  INV_X1    g0652(.A(new_n613), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT37), .B1(new_n853), .B2(new_n324), .ZN(new_n854));
  INV_X1    g0654(.A(new_n651), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n310), .A2(new_n311), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n312), .B(new_n854), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n853), .A2(new_n324), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n614), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n853), .A2(new_n651), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT100), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n330), .A2(new_n865), .A3(new_n862), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n330), .B2(new_n862), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT38), .B(new_n864), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n856), .B(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n329), .A2(new_n615), .A3(new_n616), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n861), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n869), .B(new_n859), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n869), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n423), .A2(new_n653), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n617), .A2(new_n855), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n868), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n399), .A2(new_n654), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n423), .A2(new_n426), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n887), .B1(new_n420), .B2(new_n422), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n806), .B2(new_n801), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n885), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n884), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n852), .B(new_n895), .ZN(new_n896));
  AND4_X1   g0696(.A1(new_n493), .A2(new_n576), .A3(new_n609), .A4(new_n654), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n713), .A2(new_n653), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT31), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n891), .B(new_n805), .C1(new_n897), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n802), .B1(new_n716), .B2(new_n717), .ZN(new_n906));
  NOR2_X1   g0706(.A1(KEYINPUT103), .A2(KEYINPUT40), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n906), .A2(new_n891), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n903), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n877), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n910), .A2(new_n886), .B1(new_n912), .B2(KEYINPUT40), .ZN(new_n913));
  INV_X1    g0713(.A(new_n718), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n627), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n330), .A2(new_n862), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n330), .A2(new_n865), .A3(new_n862), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n919), .B2(new_n864), .ZN(new_n920));
  INV_X1    g0720(.A(new_n868), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n905), .A2(new_n909), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n903), .B1(new_n868), .B2(new_n876), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n922), .A2(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n429), .A3(new_n718), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n915), .A2(new_n927), .A3(G330), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n896), .A2(new_n928), .B1(new_n208), .B2(new_n724), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n896), .A2(new_n928), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n849), .B1(new_n932), .B2(new_n933), .ZN(G367));
  INV_X1    g0734(.A(new_n733), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n741), .B1(new_n212), .B2(new_n371), .C1(new_n935), .C2(new_n236), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n936), .A2(new_n727), .ZN(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n343), .B1(new_n765), .B2(new_n364), .C1(new_n938), .C2(new_n815), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G97), .B2(new_n756), .ZN(new_n940));
  AOI22_X1  g0740(.A1(G303), .A2(new_n775), .B1(new_n761), .B2(G311), .ZN(new_n941));
  AOI22_X1  g0741(.A1(G283), .A2(new_n772), .B1(new_n747), .B2(G294), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n759), .A2(new_n451), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT46), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n775), .A2(G150), .B1(new_n747), .B2(G159), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n241), .B2(new_n773), .C1(new_n828), .C2(new_n762), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n755), .A2(new_n387), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n759), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(G58), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n820), .A2(G68), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n343), .B1(new_n769), .B2(G137), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n949), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n943), .A2(new_n945), .B1(new_n947), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  OR2_X1    g0756(.A1(new_n573), .A2(new_n654), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n571), .A2(new_n575), .A3(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(KEYINPUT105), .B(new_n958), .C1(new_n639), .C2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(KEYINPUT105), .B2(new_n958), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n937), .B1(new_n744), .B2(new_n956), .C1(new_n961), .C2(new_n794), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n532), .B(new_n538), .C1(new_n535), .C2(new_n654), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n509), .A2(new_n630), .A3(new_n504), .A4(new_n653), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n675), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT45), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n675), .A2(new_n965), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n660), .A3(new_n669), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n967), .A2(new_n670), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n669), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n672), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(KEYINPUT107), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n672), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n976), .B(new_n977), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n660), .A2(KEYINPUT108), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n660), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT108), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(new_n983), .A3(new_n979), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n721), .B1(new_n973), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n678), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n726), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n975), .A2(new_n965), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT42), .Z(new_n994));
  AOI21_X1  g0794(.A(new_n691), .B1(new_n965), .B2(new_n661), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n653), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n660), .A2(new_n669), .A3(new_n965), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT106), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT106), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n999), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n962), .B1(new_n992), .B2(new_n1009), .ZN(G387));
  INV_X1    g0810(.A(new_n726), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT109), .B1(new_n988), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n987), .A2(new_n1013), .A3(new_n726), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n233), .A2(G45), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT110), .Z(new_n1017));
  NOR2_X1   g0817(.A1(new_n266), .A2(G50), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n680), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT111), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n278), .B1(new_n202), .B2(new_n387), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n935), .B(new_n1017), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n731), .A2(new_n1020), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(G107), .B2(new_n212), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n741), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n727), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G303), .A2(new_n772), .B1(new_n747), .B2(G311), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n938), .B2(new_n776), .C1(new_n777), .C2(new_n762), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n950), .A2(G294), .B1(G283), .B2(new_n820), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n343), .B1(new_n763), .B2(new_n815), .C1(new_n755), .C2(new_n451), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(KEYINPUT49), .B2(new_n1036), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n348), .B1(new_n332), .B2(new_n815), .C1(new_n773), .C2(new_n202), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G97), .B2(new_n756), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n761), .A2(G159), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT112), .Z(new_n1044));
  OAI22_X1  g0844(.A1(new_n776), .A2(new_n241), .B1(new_n748), .B2(new_n266), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n371), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n820), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n950), .A2(G77), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1042), .A2(new_n1044), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n744), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1028), .B(new_n1050), .C1(new_n974), .C2(new_n739), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n679), .B1(new_n987), .B2(new_n721), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n985), .B(new_n986), .C1(new_n720), .C2(new_n702), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1015), .A2(new_n1054), .ZN(G393));
  INV_X1    g0855(.A(new_n721), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n973), .B1(new_n988), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n987), .A2(new_n971), .A3(new_n721), .A4(new_n972), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n678), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n973), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n971), .A2(KEYINPUT113), .A3(new_n972), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n1062), .A3(new_n726), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n741), .B1(new_n454), .B2(new_n212), .C1(new_n935), .C2(new_n240), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n727), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n761), .B1(new_n775), .B2(G159), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n348), .B1(new_n828), .B2(new_n815), .C1(new_n773), .C2(new_n266), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n748), .A2(new_n241), .B1(new_n765), .B2(new_n387), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n814), .B1(new_n202), .B2(new_n759), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT114), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n775), .B1(new_n761), .B2(G317), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT52), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n343), .B1(new_n815), .B2(new_n777), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n748), .A2(new_n758), .B1(new_n765), .B2(new_n451), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G294), .C2(new_n772), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n784), .B1(G283), .B2(new_n950), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1073), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1065), .B1(new_n1082), .B2(new_n740), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n965), .B2(new_n794), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1059), .A2(new_n1063), .A3(new_n1084), .ZN(G390));
  NAND3_X1  g0885(.A1(new_n906), .A2(G330), .A3(new_n891), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(KEYINPUT115), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n879), .A2(new_n882), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n893), .A2(new_n883), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n654), .B(new_n800), .C1(new_n695), .C2(new_n700), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n801), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n891), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n883), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n877), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n906), .A2(KEYINPUT115), .A3(G330), .A4(new_n891), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1089), .B1(new_n1093), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1091), .B1(new_n879), .B2(new_n882), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1088), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n850), .B(new_n626), .C1(new_n627), .C2(new_n719), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n806), .A2(new_n801), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n906), .A2(G330), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n892), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1086), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1108), .B2(new_n892), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n892), .B1(new_n719), .B2(new_n803), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1114), .A2(new_n801), .A3(new_n1086), .A4(new_n1094), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1106), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n679), .B1(new_n1105), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n738), .B1(new_n879), .B2(new_n882), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n776), .A2(new_n451), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n748), .A2(new_n364), .B1(new_n773), .B2(new_n454), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G283), .C2(new_n761), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n343), .B1(new_n765), .B2(new_n387), .C1(new_n600), .C2(new_n815), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1125), .B(new_n785), .C1(G68), .C2(new_n756), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n343), .B1(new_n769), .B2(G125), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n755), .B2(new_n241), .C1(new_n833), .C2(new_n776), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  INV_X1    g0929(.A(G137), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n762), .A2(new_n1129), .B1(new_n748), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n773), .A2(new_n1132), .B1(new_n829), .B2(new_n765), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n759), .A2(new_n332), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1124), .A2(new_n1126), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n727), .B1(new_n267), .B2(new_n811), .C1(new_n1137), .C2(new_n744), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1105), .A2(new_n1011), .B1(new_n1121), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1120), .A2(new_n1139), .ZN(G378));
  NOR2_X1   g0940(.A1(new_n627), .A2(new_n719), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n851), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT119), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G330), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n622), .A2(new_n624), .A3(new_n383), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n339), .A3(new_n855), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n339), .A2(new_n855), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n622), .A2(new_n624), .A3(new_n383), .A4(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n912), .A2(KEYINPUT40), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n905), .B(new_n909), .C1(new_n920), .C2(new_n921), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1145), .B(new_n1153), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1153), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n926), .B2(G330), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n895), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1153), .B1(new_n913), .B2(new_n1145), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n895), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n926), .A2(G330), .A3(new_n1157), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1144), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n679), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1144), .A2(new_n1164), .A3(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT120), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT120), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1144), .A2(new_n1164), .A3(new_n1170), .A4(KEYINPUT57), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n748), .A2(new_n833), .B1(new_n765), .B2(new_n332), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n761), .A2(G125), .B1(new_n772), .B2(G137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n759), .B2(new_n1132), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G128), .C2(new_n775), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n769), .A2(G124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n251), .A3(new_n277), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n756), .B2(G159), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n761), .A2(G116), .B1(new_n747), .B2(G97), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n364), .B2(new_n776), .C1(new_n371), .C2(new_n773), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G41), .B(new_n348), .C1(G283), .C2(new_n769), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1048), .A2(new_n952), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n755), .A2(new_n201), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT117), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT58), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n241), .B1(new_n291), .B2(G41), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1182), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n740), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n810), .A2(new_n241), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n727), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1153), .B2(new_n737), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1164), .B2(new_n726), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1172), .A2(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n892), .A2(new_n737), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n727), .B1(new_n811), .B2(G68), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G283), .A2(new_n775), .B1(new_n761), .B2(G294), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n364), .B2(new_n773), .C1(new_n451), .C2(new_n748), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n759), .A2(new_n454), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n343), .B1(new_n765), .B2(new_n371), .C1(new_n758), .C2(new_n815), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1205), .A2(new_n948), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT121), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(KEYINPUT121), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n348), .B1(new_n815), .B2(new_n1129), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1212), .B(new_n1187), .C1(G137), .C2(new_n775), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n762), .A2(new_n833), .B1(new_n748), .B2(new_n1132), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n773), .A2(new_n332), .B1(new_n765), .B2(new_n241), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1213), .B(new_n1216), .C1(new_n829), .C2(new_n759), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1210), .A2(new_n1211), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1203), .B1(new_n1218), .B2(new_n740), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1201), .A2(new_n726), .B1(new_n1202), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1117), .A2(new_n991), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1201), .A2(new_n1142), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(G381));
  AND3_X1   g1023(.A1(new_n1059), .A2(new_n1063), .A3(new_n1084), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n840), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1015), .A2(new_n1054), .A3(new_n796), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1225), .A2(new_n1227), .A3(G387), .A4(G381), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1120), .A2(new_n1139), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(G407));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1222), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1117), .A2(new_n1222), .A3(KEYINPUT60), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n678), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1220), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n840), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(G384), .A3(new_n1220), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n652), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1246), .A2(G2897), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1244), .B(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1172), .A2(G378), .A3(new_n1199), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1199), .A2(KEYINPUT123), .B1(new_n1165), .B2(new_n990), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1199), .A2(KEYINPUT123), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1229), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1246), .B1(new_n1249), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1235), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1244), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT63), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(new_n1224), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n796), .B1(new_n1015), .B2(new_n1054), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1226), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n990), .B1(new_n1058), .B2(new_n721), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n726), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G390), .A2(new_n1263), .A3(new_n962), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1258), .A2(new_n1260), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1260), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT124), .B1(new_n1257), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(new_n1269), .A2(new_n1254), .A3(new_n1256), .A4(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1246), .B(new_n1244), .C1(new_n1249), .C2(new_n1252), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1275), .A2(new_n1276), .B1(KEYINPUT62), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT126), .B1(new_n1277), .B2(new_n1274), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1254), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1267), .B(new_n1281), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n1271), .A2(new_n1273), .B1(new_n1280), .B2(new_n1282), .ZN(G405));
  NAND2_X1  g1083(.A1(G375), .A2(new_n1229), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1249), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1244), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(new_n1267), .ZN(G402));
endmodule


