//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AND2_X1   g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n214), .B1(new_n217), .B2(new_n220), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(G50), .B1(new_n209), .B2(G1), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT69), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n251), .A2(new_n257), .B1(new_n201), .B2(new_n253), .ZN(new_n258));
  OAI21_X1  g0058(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n260), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT8), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G58), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT67), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n269), .A2(new_n272), .A3(new_n209), .A4(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n256), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT9), .B(new_n258), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n264), .B2(new_n273), .ZN(new_n278));
  INV_X1    g0078(.A(new_n258), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n285), .A3(G274), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G222), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G223), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n293), .B1(new_n294), .B2(new_n291), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n285), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G190), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n276), .A2(new_n280), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(new_n290), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT72), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT70), .B(G200), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT72), .B1(new_n299), .B2(new_n306), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n301), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n278), .A2(new_n279), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(KEYINPUT9), .B1(G190), .B2(new_n299), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n308), .A2(new_n309), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .A4(new_n280), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n304), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n318), .B(new_n320), .C1(G179), .C2(new_n304), .ZN(new_n321));
  INV_X1    g0121(.A(G244), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n286), .B1(new_n322), .B2(new_n289), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n291), .A2(G232), .A3(new_n292), .ZN(new_n324));
  INV_X1    g0124(.A(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G107), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n324), .B(new_n330), .C1(new_n295), .C2(new_n223), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n323), .B1(new_n331), .B2(new_n298), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(KEYINPUT71), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n262), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n270), .A2(new_n335), .B1(new_n209), .B2(new_n294), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n209), .A2(G33), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n256), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n253), .A2(new_n294), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n254), .B(new_n255), .C1(G1), .C2(new_n209), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(new_n294), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT71), .B1(new_n332), .B2(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n332), .A2(new_n333), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n332), .A2(G190), .ZN(new_n350));
  INV_X1    g0150(.A(new_n344), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n351), .C1(new_n306), .C2(new_n332), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n321), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n287), .A2(new_n292), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n234), .A2(G1698), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n326), .A2(new_n354), .A3(new_n328), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n285), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n285), .A2(G238), .A3(new_n288), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n286), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT73), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n358), .A2(new_n360), .A3(new_n364), .A4(KEYINPUT13), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n356), .A2(new_n357), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n298), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n286), .A2(new_n359), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n333), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n362), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT13), .B1(new_n358), .B2(new_n360), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT14), .B1(new_n375), .B2(G169), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n377), .B(new_n319), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n372), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n342), .A2(new_n222), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n222), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n383), .A2(new_n252), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n253), .A2(new_n381), .A3(new_n382), .A4(new_n222), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n262), .A2(G50), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n222), .A2(G20), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n294), .C2(new_n338), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n389), .A2(new_n390), .A3(new_n256), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n389), .B2(new_n256), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n379), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n373), .A2(new_n364), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT73), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(G190), .A4(new_n374), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n375), .B2(G200), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND4_X1   g0200(.A1(new_n317), .A2(new_n353), .A3(new_n394), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n269), .A2(new_n272), .A3(new_n342), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n253), .B1(new_n269), .B2(new_n272), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n268), .A2(KEYINPUT67), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n270), .A2(new_n271), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n252), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n269), .A2(new_n272), .A3(new_n342), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT76), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(G58), .A2(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(G20), .B1(new_n412), .B2(new_n218), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT75), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n262), .A2(G159), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT7), .B1(new_n329), .B2(new_n209), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT7), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n420), .B(G20), .C1(new_n326), .C2(new_n328), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n275), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n418), .A2(new_n422), .A3(KEYINPUT16), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n411), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n326), .A2(new_n328), .A3(G226), .A4(G1698), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n326), .A2(new_n328), .A3(G223), .A4(new_n292), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n298), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n285), .A2(G232), .A3(new_n288), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n286), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n433), .A2(G190), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n433), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n428), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n433), .A2(G190), .A3(new_n436), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n298), .B2(new_n432), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(KEYINPUT77), .C1(new_n442), .C2(new_n438), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n427), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(G179), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n319), .B2(new_n442), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT18), .B1(new_n427), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n413), .A2(new_n415), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n420), .B1(new_n291), .B2(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n222), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n424), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n426), .A3(new_n256), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n405), .A2(new_n410), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n449), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n427), .A2(new_n444), .A3(KEYINPUT17), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n447), .A2(new_n451), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n401), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(G1698), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n326), .A2(new_n328), .A3(G244), .A4(new_n292), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n471), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n298), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n208), .B(G45), .C1(new_n281), .C2(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(KEYINPUT79), .A3(new_n208), .A4(G45), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n215), .B2(new_n284), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n481), .A2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n480), .A2(new_n483), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G257), .B(new_n285), .C1(new_n478), .C2(new_n486), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n477), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G200), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n252), .A2(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n208), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n252), .A2(new_n494), .A3(new_n255), .A4(new_n254), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n496), .B2(G97), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n335), .A2(new_n294), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n500), .A2(new_n501), .A3(G107), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n499), .B1(new_n508), .B2(G20), .ZN(new_n509));
  OAI21_X1  g0309(.A(G107), .B1(new_n419), .B2(new_n421), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n498), .B1(new_n511), .B2(new_n256), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n477), .A2(new_n490), .A3(G190), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n492), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n491), .A2(new_n319), .ZN(new_n515));
  INV_X1    g0315(.A(new_n499), .ZN(new_n516));
  XNOR2_X1  g0316(.A(G97), .B(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n506), .B1(new_n517), .B2(new_n500), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(new_n209), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n502), .B1(new_n456), .B2(new_n457), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n256), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n497), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n477), .A2(new_n490), .A3(new_n333), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n515), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n326), .A2(new_n328), .A3(G244), .A4(G1698), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n326), .A2(new_n328), .A3(G238), .A4(new_n292), .ZN(new_n527));
  INV_X1    g0327(.A(G116), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n325), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n298), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n225), .B1(new_n282), .B2(G1), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n208), .A2(new_n484), .A3(G45), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n285), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n307), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n209), .B1(new_n357), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n504), .A2(new_n224), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n326), .A2(new_n328), .A3(new_n209), .A4(G68), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n538), .B1(new_n338), .B2(new_n501), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n256), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n337), .A2(new_n253), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n496), .A2(G87), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n535), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n531), .B2(new_n298), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n537), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n337), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n496), .A2(KEYINPUT80), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n495), .B2(new_n337), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n545), .A2(new_n554), .A3(new_n546), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n333), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(G169), .C2(new_n550), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n525), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n326), .A2(new_n328), .A3(new_n209), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n291), .A2(new_n564), .A3(new_n209), .A4(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n209), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n502), .A2(KEYINPUT23), .A3(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n529), .A2(new_n209), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT82), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n572), .B1(new_n563), .B2(new_n565), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT24), .B1(new_n578), .B2(KEYINPUT82), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n573), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n577), .B(new_n256), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT25), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n252), .B2(G107), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n252), .A2(new_n582), .A3(G107), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n584), .A2(new_n585), .B1(new_n502), .B2(new_n495), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(G1698), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n326), .A2(new_n328), .A3(G250), .A4(new_n292), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n298), .ZN(new_n593));
  OAI211_X1 g0393(.A(G264), .B(new_n285), .C1(new_n478), .C2(new_n486), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n488), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n319), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G179), .B2(new_n595), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n588), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n275), .B1(new_n600), .B2(new_n576), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n574), .A2(new_n575), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(KEYINPUT24), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n586), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT83), .B1(new_n595), .B2(G190), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n595), .A2(new_n438), .ZN(new_n607));
  INV_X1    g0407(.A(new_n594), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n298), .B2(new_n592), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT83), .ZN(new_n610));
  INV_X1    g0410(.A(G190), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n488), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n599), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n528), .A2(G20), .ZN(new_n616));
  INV_X1    g0416(.A(G13), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n616), .A2(G1), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n471), .B(new_n209), .C1(G33), .C2(new_n501), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n256), .A3(new_n616), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(KEYINPUT20), .A3(new_n256), .A4(new_n616), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n496), .A2(KEYINPUT81), .A3(G116), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT81), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n495), .B2(new_n528), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n326), .A2(new_n328), .A3(G264), .A4(G1698), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n326), .A2(new_n328), .A3(G257), .A4(new_n292), .ZN(new_n631));
  INV_X1    g0431(.A(G303), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n291), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n298), .ZN(new_n634));
  OAI211_X1 g0434(.A(G270), .B(new_n285), .C1(new_n478), .C2(new_n486), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n488), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n629), .A2(new_n636), .A3(KEYINPUT21), .A4(G169), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n488), .A2(new_n635), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n629), .A2(G179), .A3(new_n634), .A4(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n629), .B1(G200), .B2(new_n636), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n611), .B2(new_n636), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n629), .A2(G169), .A3(new_n636), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT21), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n561), .A2(new_n615), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n470), .A2(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n321), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n317), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n316), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n450), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n463), .B1(new_n462), .B2(new_n449), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n427), .A2(new_n444), .A3(KEYINPUT17), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT17), .B1(new_n427), .B2(new_n444), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n349), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(new_n400), .B1(new_n379), .B2(new_n393), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n656), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n649), .B1(new_n653), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n515), .A2(new_n523), .A3(new_n522), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT84), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n536), .A2(new_n667), .A3(new_n307), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT84), .B1(new_n550), .B2(new_n306), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n551), .A4(new_n548), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n665), .A2(new_n666), .A3(new_n559), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n552), .A2(new_n559), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n672), .B2(new_n524), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n559), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n640), .A2(new_n645), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT85), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n605), .A2(new_n676), .A3(new_n597), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT85), .B1(new_n588), .B2(new_n598), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n670), .A2(new_n559), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n525), .A2(new_n614), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n674), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n664), .B1(new_n469), .B2(new_n683), .ZN(G369));
  NAND3_X1  g0484(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n605), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n615), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT88), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n599), .A2(new_n690), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n615), .A2(new_n691), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT88), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n629), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT87), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n675), .A2(new_n642), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n675), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n640), .A2(new_n645), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n690), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n696), .B2(new_n698), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n677), .A2(new_n678), .A3(new_n701), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0515(.A(new_n212), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n540), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n220), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n593), .A2(new_n594), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n536), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n638), .A2(G179), .A3(new_n634), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n477), .A2(new_n490), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n609), .A2(KEYINPUT90), .A3(new_n550), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n491), .A2(new_n595), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT93), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n636), .A2(new_n333), .A3(new_n536), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n731), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT91), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n491), .A2(new_n636), .A3(new_n333), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(KEYINPUT91), .A3(new_n728), .A4(new_n725), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT92), .B(KEYINPUT30), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n561), .A2(new_n615), .A3(new_n646), .A4(new_n701), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT94), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n742), .B1(new_n729), .B2(new_n738), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(KEYINPUT94), .A3(new_n741), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n690), .B1(new_n753), .B2(new_n737), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n746), .B(new_n748), .C1(new_n754), .C2(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n673), .A2(new_n559), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n599), .A2(new_n676), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n588), .A2(new_n598), .A3(KEYINPUT85), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n709), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n680), .B1(new_n605), .B2(new_n613), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n525), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n671), .B(new_n757), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n690), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n599), .A2(new_n645), .A3(new_n640), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n514), .A2(new_n524), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT96), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n514), .A2(new_n524), .A3(KEYINPUT96), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n767), .A2(new_n761), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT26), .B1(new_n680), .B2(new_n524), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n560), .A2(new_n665), .A3(new_n666), .ZN(new_n774));
  AND3_X1   g0574(.A1(new_n773), .A2(new_n774), .A3(new_n559), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n701), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT29), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n766), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n756), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n722), .B1(new_n779), .B2(G1), .ZN(G364));
  INV_X1    g0580(.A(new_n706), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n617), .A2(G20), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n208), .B1(new_n782), .B2(G45), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n717), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G330), .B2(new_n705), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n212), .A2(new_n291), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n788), .A2(new_n206), .B1(G116), .B2(new_n212), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n245), .A2(G45), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n716), .A2(new_n291), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n220), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n282), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n789), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n209), .B1(KEYINPUT97), .B2(new_n319), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n319), .A2(KEYINPUT97), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n255), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT98), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n785), .B1(new_n795), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n209), .A2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n306), .A2(new_n806), .A3(G179), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT102), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT102), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G107), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G179), .A2(G200), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n209), .B1(new_n814), .B2(G190), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n501), .ZN(new_n816));
  NAND3_X1  g0616(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G190), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n611), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n819), .A2(new_n222), .B1(new_n821), .B2(new_n201), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n805), .A2(new_n814), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT100), .B(G159), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n816), .B(new_n822), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n209), .A2(new_n611), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n829), .A2(new_n306), .A3(G179), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G87), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n825), .A2(new_n826), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n333), .A2(G200), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n291), .B1(new_n834), .B2(new_n202), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n805), .A2(new_n833), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n832), .B(new_n835), .C1(new_n842), .C2(G77), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n813), .A2(new_n827), .A3(new_n831), .A4(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n811), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(G311), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT33), .B(G317), .Z(new_n848));
  INV_X1    g0648(.A(G326), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n819), .A2(new_n848), .B1(new_n821), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n815), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(G294), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(G329), .ZN(new_n853));
  INV_X1    g0653(.A(G322), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n329), .B1(new_n823), .B2(new_n853), .C1(new_n834), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G303), .B2(new_n830), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n847), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n844), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n804), .B1(new_n858), .B2(new_n798), .ZN(new_n859));
  INV_X1    g0659(.A(new_n801), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n705), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n787), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G396));
  NAND2_X1  g0663(.A1(new_n812), .A2(G87), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n821), .A2(new_n632), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n816), .B(new_n865), .C1(G283), .C2(new_n818), .ZN(new_n866));
  INV_X1    g0666(.A(G311), .ZN(new_n867));
  INV_X1    g0667(.A(G294), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n329), .B1(new_n823), .B2(new_n867), .C1(new_n834), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n830), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(new_n502), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n869), .B(new_n871), .C1(G116), .C2(new_n842), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n874));
  INV_X1    g0674(.A(new_n834), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(G143), .B1(G137), .B2(new_n820), .ZN(new_n876));
  INV_X1    g0676(.A(G150), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n876), .B1(new_n877), .B2(new_n819), .C1(new_n841), .C2(new_n824), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT34), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(KEYINPUT34), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n812), .A2(G68), .ZN(new_n882));
  INV_X1    g0682(.A(G132), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n291), .B1(new_n815), .B2(new_n202), .C1(new_n883), .C2(new_n823), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(G50), .B2(new_n830), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n874), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n798), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n798), .A2(new_n799), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n889), .B(new_n785), .C1(G77), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n701), .A2(new_n344), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n348), .A2(new_n345), .B1(new_n352), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n345), .A2(new_n348), .A3(new_n690), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT104), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n352), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n349), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT104), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n345), .A2(new_n348), .A3(new_n690), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n799), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n764), .A2(new_n903), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n896), .A2(new_n690), .A3(new_n901), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n683), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(new_n756), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n785), .B1(new_n907), .B2(new_n756), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(G384));
  NOR2_X1   g0711(.A1(new_n782), .A2(new_n208), .ZN(new_n912));
  INV_X1    g0712(.A(G330), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n408), .A2(new_n409), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n460), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n689), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n659), .B2(new_n656), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n462), .B1(new_n449), .B2(new_n689), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n445), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n449), .B2(new_n689), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n445), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n915), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT107), .ZN(new_n927));
  INV_X1    g0727(.A(new_n918), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n466), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n445), .A2(new_n920), .A3(new_n921), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n445), .A2(new_n923), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n921), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(KEYINPUT38), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n926), .A2(new_n927), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n927), .B1(new_n926), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND4_X1   g0736(.A1(KEYINPUT94), .A2(new_n739), .A3(new_n741), .A4(new_n743), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT94), .B1(new_n751), .B2(new_n741), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n737), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n748), .C1(new_n754), .C2(KEYINPUT31), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n701), .A2(new_n393), .ZN(new_n942));
  OAI21_X1  g0742(.A(G169), .B1(new_n370), .B2(new_n396), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n377), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n375), .A2(KEYINPUT14), .A3(G169), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n944), .A2(new_n945), .B1(new_n366), .B2(new_n371), .ZN(new_n946));
  INV_X1    g0746(.A(new_n393), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n400), .B(new_n942), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n942), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n398), .A2(new_n399), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n379), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT105), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT106), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT105), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n394), .A2(new_n954), .A3(new_n400), .A4(new_n942), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n953), .B1(new_n952), .B2(new_n955), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n941), .A2(new_n959), .A3(new_n902), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n914), .B1(new_n936), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n427), .A2(new_n688), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n659), .B2(new_n656), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n921), .B1(new_n445), .B2(new_n920), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n922), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n915), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n914), .B1(new_n967), .B2(new_n933), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n968), .A2(new_n941), .A3(new_n902), .A4(new_n959), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT31), .B1(new_n939), .B2(new_n701), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n701), .A2(KEYINPUT31), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n753), .B2(new_n737), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n972), .A2(new_n974), .A3(new_n747), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n469), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n913), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n971), .B2(new_n976), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n919), .A2(new_n925), .A3(new_n915), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT38), .B1(new_n929), .B2(new_n932), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT107), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n926), .A2(new_n927), .A3(new_n933), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n900), .B1(new_n683), .B2(new_n906), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n984), .A3(new_n959), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT39), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n466), .A2(new_n962), .ZN(new_n987));
  INV_X1    g0787(.A(new_n965), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n930), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT38), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n979), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n379), .A2(new_n393), .A3(new_n690), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT108), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n688), .B1(new_n654), .B2(new_n655), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n985), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n664), .B1(new_n778), .B2(new_n469), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n997), .B(new_n998), .Z(new_n999));
  AOI21_X1  g0799(.A(new_n912), .B1(new_n978), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n999), .B2(new_n978), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n528), .A4(new_n217), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT36), .Z(new_n1005));
  OR3_X1    g0805(.A1(new_n220), .A2(new_n294), .A3(new_n412), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n201), .A2(G68), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(G1), .A3(new_n617), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1001), .A2(new_n1005), .A3(new_n1009), .ZN(G367));
  OAI22_X1  g0810(.A1(new_n841), .A2(new_n201), .B1(new_n294), .B2(new_n808), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n851), .A2(G68), .B1(G143), .B2(new_n820), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n824), .B2(new_n819), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n870), .A2(new_n202), .ZN(new_n1014));
  INV_X1    g0814(.A(G137), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n291), .B1(new_n823), .B2(new_n1015), .C1(new_n834), .C2(new_n877), .ZN(new_n1016));
  NOR4_X1   g0816(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT113), .Z(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n329), .B1(new_n823), .B2(new_n1019), .C1(new_n834), .C2(new_n632), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n808), .A2(new_n501), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G283), .C2(new_n842), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n851), .A2(G107), .B1(G311), .B2(new_n820), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n868), .B2(new_n819), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n870), .A2(new_n528), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(KEYINPUT46), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1026), .C1(KEYINPUT46), .C2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1018), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT47), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n798), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n548), .A2(new_n690), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n681), .A2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n559), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n801), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n803), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n791), .A2(new_n240), .B1(new_n716), .B2(new_n553), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n717), .B(new_n784), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1030), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n710), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n699), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n711), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(new_n706), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n779), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT45), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n699), .A2(new_n1040), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n712), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n524), .A2(new_n690), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n770), .B(new_n771), .C1(new_n512), .C2(new_n690), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1046), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n1053), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1049), .A2(KEYINPUT44), .A3(new_n1054), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT44), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n713), .B2(new_n1053), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n707), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1057), .A2(new_n1061), .A3(new_n708), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1045), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT112), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1064), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n708), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT112), .B1(new_n1070), .B2(new_n1045), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n779), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n717), .B(KEYINPUT41), .Z(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n784), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT43), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n1078));
  NAND3_X1  g0878(.A1(new_n1033), .A2(new_n1034), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1053), .A2(new_n588), .A3(new_n598), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n701), .B1(new_n1081), .B2(new_n524), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n711), .A2(new_n1053), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT42), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT42), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  MUX2_X1   g0887(.A(new_n1080), .B(new_n1079), .S(new_n1087), .Z(new_n1088));
  NAND2_X1  g0888(.A1(new_n707), .A2(new_n1053), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1039), .B1(new_n1075), .B2(new_n1091), .ZN(G387));
  NAND2_X1  g0892(.A1(new_n1043), .A2(new_n784), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT114), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n788), .A2(new_n719), .B1(G107), .B2(new_n212), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n237), .A2(new_n282), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n719), .ZN(new_n1097));
  AOI211_X1 g0897(.A(G45), .B(new_n1097), .C1(G68), .C2(G77), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n270), .A2(G50), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT50), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n792), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1095), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(G159), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n291), .B1(new_n821), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n842), .B2(G68), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n406), .A2(new_n407), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n818), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(new_n811), .C2(new_n501), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n851), .A2(new_n553), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n201), .B2(new_n834), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT116), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n830), .A2(G77), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n877), .B2(new_n823), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1108), .A2(new_n1111), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n329), .B1(new_n823), .B2(new_n849), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n875), .A2(G317), .B1(G311), .B2(new_n818), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n854), .B2(new_n821), .C1(new_n841), .C2(new_n632), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT48), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n830), .A2(G294), .B1(G283), .B2(new_n851), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT49), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1117), .B(new_n1126), .C1(G116), .C2(new_n807), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1116), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n798), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n785), .B1(new_n803), .B2(new_n1102), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT117), .Z(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n700), .B2(new_n801), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1094), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1045), .A2(new_n718), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n779), .B2(new_n1043), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(G393));
  NAND2_X1  g0937(.A1(new_n791), .A2(new_n248), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n501), .B2(new_n212), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n785), .B1(new_n1139), .B2(new_n803), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n821), .A2(new_n877), .B1(new_n834), .B2(new_n1103), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT51), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n815), .A2(new_n294), .ZN(new_n1143));
  INV_X1    g0943(.A(G143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n291), .B1(new_n823), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G50), .C2(new_n818), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n842), .A2(new_n268), .B1(G68), .B2(new_n830), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n864), .A2(new_n1142), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n329), .B1(new_n823), .B2(new_n854), .C1(new_n819), .C2(new_n632), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G116), .B2(new_n851), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n842), .A2(G294), .B1(G283), .B2(new_n830), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n813), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n875), .A2(G311), .B1(G317), .B2(new_n820), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT52), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1140), .B1(new_n1155), .B2(new_n798), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1053), .B2(new_n860), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1070), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n783), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1070), .A2(KEYINPUT112), .A3(new_n1045), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n718), .B1(new_n1158), .B2(new_n1044), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1159), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G390));
  NAND2_X1  g0965(.A1(new_n991), .A2(new_n994), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n952), .A2(new_n955), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT106), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n984), .A2(new_n1168), .A3(new_n956), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n993), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT118), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n993), .B1(new_n967), .B2(new_n933), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1168), .A2(new_n956), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n895), .B1(new_n776), .B2(new_n902), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n755), .A2(new_n959), .A3(G330), .A4(new_n902), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1172), .A2(new_n1173), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n941), .A2(new_n959), .A3(G330), .A4(new_n902), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n991), .A2(new_n994), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1170), .B1(new_n979), .B2(new_n990), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1181), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n776), .A2(new_n902), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n959), .B1(new_n1188), .B2(new_n895), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1166), .A2(new_n1171), .B1(new_n1189), .B2(new_n1174), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1173), .B1(new_n1190), .B2(new_n1178), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1166), .A2(new_n799), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n785), .B1(new_n891), .B2(new_n1106), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n821), .A2(new_n845), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1143), .B(new_n1195), .C1(G107), .C2(new_n818), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n842), .A2(G97), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n329), .B1(new_n823), .B2(new_n868), .C1(new_n834), .C2(new_n528), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G87), .B2(new_n830), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n882), .A2(new_n1196), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n830), .A2(G150), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT53), .ZN(new_n1202));
  INV_X1    g1002(.A(G128), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n821), .A2(new_n1203), .B1(new_n815), .B2(new_n1103), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G137), .B2(new_n818), .ZN(new_n1205));
  INV_X1    g1005(.A(G125), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n291), .B1(new_n823), .B2(new_n1206), .C1(new_n834), .C2(new_n883), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT54), .B(G143), .Z(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n842), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1205), .B(new_n1209), .C1(new_n201), .C2(new_n808), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1200), .B1(new_n1202), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1194), .B1(new_n1211), .B2(new_n798), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1192), .A2(new_n784), .B1(new_n1193), .B2(new_n1212), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT39), .B1(new_n967), .B2(new_n933), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n993), .B1(new_n959), .B2(new_n984), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1177), .B(new_n1178), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT118), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n1186), .A3(new_n1179), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n470), .A2(new_n766), .A3(new_n777), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n941), .A2(G330), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n664), .C1(new_n1222), .C2(new_n469), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n939), .A2(new_n701), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT31), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n747), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n913), .B1(new_n1227), .B2(new_n940), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n959), .B1(new_n1228), .B2(new_n902), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1178), .A2(new_n1176), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n984), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n755), .A2(G330), .A3(new_n902), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1175), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1180), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1224), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n718), .B1(new_n1220), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT119), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1180), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n984), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1175), .B1(new_n1222), .B2(new_n903), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1223), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1219), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1237), .A2(new_n1238), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1238), .B1(new_n1237), .B2(new_n1245), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1213), .B1(new_n1246), .B2(new_n1247), .ZN(G378));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n651), .A2(new_n321), .A3(new_n652), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n312), .A2(new_n688), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1251), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n651), .A2(new_n321), .A3(new_n652), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1255), .B(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1168), .A2(new_n902), .A3(new_n956), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n975), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT40), .B1(new_n1259), .B2(new_n983), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n969), .A2(G330), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n913), .B1(new_n1259), .B2(new_n968), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1256), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1255), .B(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n961), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1262), .A2(new_n1266), .A3(new_n997), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n997), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT57), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1223), .B(KEYINPUT122), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1192), .B2(new_n1243), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1249), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1223), .B(KEYINPUT122), .Z(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1220), .B2(new_n1236), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n997), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1262), .A2(new_n1266), .A3(new_n997), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1279), .A3(KEYINPUT123), .A4(KEYINPUT57), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1245), .A2(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n717), .B1(new_n1282), .B2(KEYINPUT57), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1279), .A2(new_n784), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n784), .B(new_n717), .C1(new_n201), .C2(new_n890), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n291), .A2(G41), .ZN(new_n1287));
  AOI211_X1 g1087(.A(G50), .B(new_n1287), .C1(new_n325), .C2(new_n281), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n842), .A2(G137), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n875), .A2(G128), .B1(new_n851), .B2(G150), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(G125), .A2(new_n820), .B1(new_n818), .B2(G132), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n830), .A2(new_n1208), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT59), .ZN(new_n1294));
  INV_X1    g1094(.A(G124), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n823), .A2(new_n1295), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(G33), .A3(G41), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1294), .B(new_n1297), .C1(new_n808), .C2(new_n824), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1293), .A2(KEYINPUT59), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT58), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1112), .A2(new_n1287), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1301), .A2(KEYINPUT120), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n842), .A2(new_n553), .B1(G58), .B2(new_n807), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n834), .A2(new_n502), .B1(new_n823), .B2(new_n845), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n819), .A2(new_n501), .B1(new_n821), .B2(new_n528), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1304), .B(new_n1305), .C1(G68), .C2(new_n851), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1301), .A2(KEYINPUT120), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1302), .A2(new_n1303), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1298), .A2(new_n1299), .B1(new_n1300), .B2(new_n1308), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1288), .B(new_n1309), .C1(new_n1300), .C2(new_n1308), .ZN(new_n1310));
  OAI221_X1 g1110(.A(new_n1286), .B1(new_n1130), .B2(new_n1310), .C1(new_n1265), .C2(new_n800), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(KEYINPUT121), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1285), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1284), .A2(new_n1314), .ZN(G375));
  NOR2_X1   g1115(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1223), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1318), .A2(new_n1243), .A3(new_n1073), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n785), .B1(new_n891), .B2(G68), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n329), .B1(new_n823), .B2(new_n632), .C1(new_n834), .C2(new_n845), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n842), .B2(G107), .ZN(new_n1322));
  OAI221_X1 g1122(.A(new_n1109), .B1(new_n821), .B2(new_n868), .C1(new_n528), .C2(new_n819), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1322), .B(new_n1324), .C1(new_n501), .C2(new_n870), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n811), .A2(new_n294), .ZN(new_n1326));
  OAI221_X1 g1126(.A(new_n291), .B1(new_n823), .B2(new_n1203), .C1(new_n834), .C2(new_n1015), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(G58), .B2(new_n807), .ZN(new_n1328));
  OAI221_X1 g1128(.A(new_n1328), .B1(new_n877), .B2(new_n841), .C1(new_n1103), .C2(new_n870), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1208), .A2(new_n818), .ZN(new_n1330));
  OAI221_X1 g1130(.A(new_n1330), .B1(new_n201), .B2(new_n815), .C1(new_n821), .C2(new_n883), .ZN(new_n1331));
  OAI22_X1  g1131(.A1(new_n1325), .A2(new_n1326), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1320), .B1(new_n1332), .B2(new_n798), .ZN(new_n1333));
  XOR2_X1   g1133(.A(new_n1333), .B(KEYINPUT124), .Z(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n959), .B2(new_n800), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1335), .B1(new_n1316), .B2(new_n783), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1319), .A2(new_n1336), .ZN(G381));
  NAND2_X1  g1137(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1338), .A2(new_n1213), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(G375), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1134), .A2(new_n862), .A3(new_n1136), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(new_n1164), .A3(new_n910), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(G387), .A2(G381), .A3(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1342), .B1(KEYINPUT125), .B2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1347), .B1(KEYINPUT125), .B2(new_n1346), .ZN(G407));
  OAI211_X1 g1148(.A(G407), .B(G213), .C1(G343), .C2(new_n1342), .ZN(G409));
  AOI21_X1  g1149(.A(new_n862), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1344), .A2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1039), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n779), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n783), .B1(new_n1355), .B2(new_n1073), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1353), .B1(new_n1356), .B2(new_n1090), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1357), .A2(G390), .ZN(new_n1358));
  AOI211_X1 g1158(.A(new_n1353), .B(new_n1164), .C1(new_n1356), .C2(new_n1090), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1352), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G387), .A2(new_n1164), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1357), .A2(G390), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1361), .A2(new_n1351), .A3(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1360), .A2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(G213), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1365), .A2(G343), .ZN(new_n1366));
  OAI211_X1 g1166(.A(G378), .B(new_n1314), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1367));
  AND2_X1   g1167(.A1(new_n1282), .A2(new_n1074), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1339), .B1(new_n1368), .B2(new_n1313), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1366), .B1(new_n1367), .B2(new_n1369), .ZN(new_n1370));
  AND2_X1   g1170(.A1(new_n1236), .A2(KEYINPUT60), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n718), .B1(new_n1371), .B2(new_n1318), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1236), .A2(KEYINPUT60), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1373), .A2(new_n1317), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1336), .B1(new_n1372), .B2(new_n1374), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1375), .A2(G384), .ZN(new_n1376));
  AOI211_X1 g1176(.A(new_n910), .B(new_n1336), .C1(new_n1372), .C2(new_n1374), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  AND2_X1   g1178(.A1(new_n1370), .A2(new_n1378), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1364), .B1(KEYINPUT63), .B2(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT126), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1382));
  INV_X1    g1182(.A(new_n1366), .ZN(new_n1383));
  AND4_X1   g1183(.A1(new_n1381), .A2(new_n1382), .A3(new_n1378), .A4(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1184(.A(new_n1381), .B1(new_n1370), .B2(new_n1378), .ZN(new_n1385));
  OR3_X1    g1185(.A1(new_n1384), .A2(new_n1385), .A3(KEYINPUT63), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT61), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1366), .A2(G2897), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1388), .ZN(new_n1389));
  OAI21_X1  g1189(.A(new_n1389), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n717), .B1(new_n1373), .B2(new_n1317), .ZN(new_n1391));
  AOI21_X1  g1191(.A(new_n1391), .B1(new_n1317), .B2(new_n1373), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n910), .B1(new_n1392), .B2(new_n1336), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1375), .A2(G384), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1393), .A2(new_n1394), .A3(new_n1388), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1390), .A2(new_n1395), .ZN(new_n1396));
  OAI21_X1  g1196(.A(new_n1387), .B1(new_n1396), .B2(new_n1370), .ZN(new_n1397));
  INV_X1    g1197(.A(new_n1397), .ZN(new_n1398));
  NAND3_X1  g1198(.A1(new_n1380), .A2(new_n1386), .A3(new_n1398), .ZN(new_n1399));
  INV_X1    g1199(.A(KEYINPUT62), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1400), .B1(new_n1384), .B2(new_n1385), .ZN(new_n1401));
  AOI21_X1  g1201(.A(new_n1400), .B1(new_n1370), .B2(new_n1378), .ZN(new_n1402));
  NOR2_X1   g1202(.A1(new_n1397), .A2(new_n1402), .ZN(new_n1403));
  NAND3_X1  g1203(.A1(new_n1401), .A2(KEYINPUT127), .A3(new_n1403), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1404), .A2(new_n1364), .ZN(new_n1405));
  AOI21_X1  g1205(.A(KEYINPUT127), .B1(new_n1401), .B2(new_n1403), .ZN(new_n1406));
  OAI21_X1  g1206(.A(new_n1399), .B1(new_n1405), .B2(new_n1406), .ZN(G405));
  NAND2_X1  g1207(.A1(G375), .A2(new_n1339), .ZN(new_n1408));
  NAND2_X1  g1208(.A1(new_n1408), .A2(new_n1367), .ZN(new_n1409));
  OR2_X1    g1209(.A1(new_n1409), .A2(new_n1378), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1409), .A2(new_n1378), .ZN(new_n1411));
  NAND2_X1  g1211(.A1(new_n1410), .A2(new_n1411), .ZN(new_n1412));
  XNOR2_X1  g1212(.A(new_n1412), .B(new_n1364), .ZN(G402));
endmodule


