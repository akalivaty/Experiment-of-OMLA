

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771;

  XNOR2_X1 U374 ( .A(KEYINPUT85), .B(KEYINPUT46), .ZN(n350) );
  NOR2_X2 U375 ( .A1(n615), .A2(n434), .ZN(n367) );
  XNOR2_X2 U376 ( .A(n479), .B(n478), .ZN(n730) );
  OR2_X2 U377 ( .A1(n594), .A2(n713), .ZN(n587) );
  INV_X1 U378 ( .A(n689), .ZN(n422) );
  NAND2_X1 U379 ( .A1(n552), .A2(n550), .ZN(n689) );
  NAND2_X1 U380 ( .A1(n623), .A2(n646), .ZN(n734) );
  XNOR2_X1 U381 ( .A(n409), .B(n350), .ZN(n412) );
  INV_X1 U382 ( .A(n657), .ZN(n568) );
  NAND2_X1 U383 ( .A1(n656), .A2(n647), .ZN(n409) );
  XNOR2_X1 U384 ( .A(n433), .B(KEYINPUT39), .ZN(n609) );
  NAND2_X1 U385 ( .A1(n408), .A2(n608), .ZN(n433) );
  XNOR2_X1 U386 ( .A(n581), .B(n580), .ZN(n582) );
  NOR2_X1 U387 ( .A1(n579), .A2(n593), .ZN(n581) );
  XNOR2_X1 U388 ( .A(n546), .B(KEYINPUT105), .ZN(n594) );
  XNOR2_X1 U389 ( .A(n534), .B(G137), .ZN(n761) );
  XNOR2_X1 U390 ( .A(KEYINPUT91), .B(KEYINPUT17), .ZN(n484) );
  INV_X2 U391 ( .A(G953), .ZN(n505) );
  AND2_X1 U392 ( .A1(n733), .A2(n573), .ZN(n436) );
  NAND2_X1 U393 ( .A1(n353), .A2(n626), .ZN(n627) );
  INV_X1 U394 ( .A(n734), .ZN(n757) );
  NAND2_X1 U395 ( .A1(n403), .A2(n410), .ZN(n411) );
  AND2_X1 U396 ( .A1(n382), .A2(n384), .ZN(n366) );
  NOR2_X1 U397 ( .A1(n352), .A2(n622), .ZN(n351) );
  AND2_X1 U398 ( .A1(n380), .A2(n377), .ZN(n376) );
  AND2_X1 U399 ( .A1(n602), .A2(n601), .ZN(n407) );
  XNOR2_X1 U400 ( .A(n563), .B(n562), .ZN(n655) );
  INV_X1 U401 ( .A(n609), .ZN(n354) );
  NAND2_X1 U402 ( .A1(n609), .A2(n422), .ZN(n402) );
  XNOR2_X1 U403 ( .A(n614), .B(n613), .ZN(n647) );
  AND2_X1 U404 ( .A1(n595), .A2(n544), .ZN(n612) );
  XNOR2_X1 U405 ( .A(n604), .B(n603), .ZN(n712) );
  NAND2_X1 U406 ( .A1(n604), .A2(n610), .ZN(n583) );
  NAND2_X2 U407 ( .A1(n371), .A2(n370), .ZN(n604) );
  AND2_X1 U408 ( .A1(n372), .A2(n375), .ZN(n371) );
  BUF_X1 U409 ( .A(n543), .Z(n544) );
  OR2_X1 U410 ( .A1(n651), .A2(G902), .ZN(n460) );
  XNOR2_X1 U411 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U412 ( .A(n487), .B(G134), .ZN(n534) );
  NAND2_X1 U413 ( .A1(n621), .A2(KEYINPUT2), .ZN(n622) );
  XNOR2_X1 U414 ( .A(KEYINPUT78), .B(KEYINPUT89), .ZN(n481) );
  XNOR2_X1 U415 ( .A(G131), .B(KEYINPUT74), .ZN(n414) );
  NAND2_X1 U416 ( .A1(n623), .A2(n351), .ZN(n353) );
  INV_X1 U417 ( .A(n646), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n355), .B(KEYINPUT28), .ZN(n595) );
  NOR2_X1 U419 ( .A1(n594), .A2(n593), .ZN(n355) );
  INV_X1 U420 ( .A(n424), .ZN(n356) );
  BUF_X1 U421 ( .A(n679), .Z(n357) );
  XNOR2_X1 U422 ( .A(n572), .B(n425), .ZN(n742) );
  XNOR2_X1 U423 ( .A(n426), .B(KEYINPUT102), .ZN(n679) );
  NOR2_X1 U424 ( .A1(n555), .A2(n588), .ZN(n545) );
  XNOR2_X2 U425 ( .A(n411), .B(n620), .ZN(n623) );
  XNOR2_X1 U426 ( .A(n546), .B(KEYINPUT6), .ZN(n579) );
  XNOR2_X2 U427 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n369) );
  XNOR2_X2 U428 ( .A(G146), .B(G125), .ZN(n488) );
  XNOR2_X1 U429 ( .A(n599), .B(KEYINPUT83), .ZN(n406) );
  INV_X1 U430 ( .A(n649), .ZN(n379) );
  NOR2_X1 U431 ( .A1(n542), .A2(KEYINPUT44), .ZN(n378) );
  NAND2_X1 U432 ( .A1(n650), .A2(n435), .ZN(n404) );
  XNOR2_X1 U433 ( .A(G119), .B(G116), .ZN(n467) );
  XNOR2_X1 U434 ( .A(n488), .B(KEYINPUT10), .ZN(n516) );
  XNOR2_X1 U435 ( .A(n394), .B(n393), .ZN(n529) );
  INV_X1 U436 ( .A(KEYINPUT8), .ZN(n393) );
  NAND2_X1 U437 ( .A1(n422), .A2(n584), .ZN(n420) );
  XNOR2_X1 U438 ( .A(G116), .B(G107), .ZN(n527) );
  INV_X1 U439 ( .A(KEYINPUT65), .ZN(n631) );
  INV_X1 U440 ( .A(KEYINPUT43), .ZN(n387) );
  AND2_X1 U441 ( .A1(n617), .A2(n616), .ZN(n388) );
  NAND2_X1 U442 ( .A1(n374), .A2(n497), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n585), .B(KEYINPUT30), .ZN(n586) );
  XNOR2_X1 U444 ( .A(n401), .B(n363), .ZN(n567) );
  XOR2_X1 U445 ( .A(n642), .B(KEYINPUT59), .Z(n643) );
  NOR2_X1 U446 ( .A1(n379), .A2(n378), .ZN(n377) );
  AND2_X1 U447 ( .A1(n578), .A2(n694), .ZN(n697) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n519) );
  XNOR2_X1 U449 ( .A(G113), .B(G143), .ZN(n517) );
  XNOR2_X1 U450 ( .A(G131), .B(G140), .ZN(n515) );
  XNOR2_X1 U451 ( .A(KEYINPUT18), .B(KEYINPUT77), .ZN(n482) );
  NAND2_X1 U452 ( .A1(n413), .A2(n412), .ZN(n410) );
  AND2_X1 U453 ( .A1(n556), .A2(n697), .ZN(n476) );
  INV_X1 U454 ( .A(n501), .ZN(n374) );
  INV_X1 U455 ( .A(G902), .ZN(n535) );
  NAND2_X1 U456 ( .A1(n544), .A2(n697), .ZN(n588) );
  XNOR2_X1 U457 ( .A(n369), .B(n399), .ZN(n465) );
  XNOR2_X1 U458 ( .A(G101), .B(KEYINPUT67), .ZN(n399) );
  XNOR2_X1 U459 ( .A(G113), .B(KEYINPUT69), .ZN(n466) );
  XNOR2_X1 U460 ( .A(n400), .B(n437), .ZN(n748) );
  INV_X1 U461 ( .A(G104), .ZN(n437) );
  XNOR2_X1 U462 ( .A(G110), .B(G107), .ZN(n400) );
  XNOR2_X1 U463 ( .A(G119), .B(G110), .ZN(n451) );
  XNOR2_X1 U464 ( .A(n465), .B(n748), .ZN(n480) );
  XOR2_X1 U465 ( .A(G131), .B(G140), .Z(n438) );
  NOR2_X1 U466 ( .A1(n420), .A2(KEYINPUT36), .ZN(n417) );
  AND2_X1 U467 ( .A1(n416), .A2(n421), .ZN(n391) );
  AND2_X1 U468 ( .A1(n419), .A2(n698), .ZN(n416) );
  NAND2_X1 U469 ( .A1(n420), .A2(KEYINPUT36), .ZN(n419) );
  XNOR2_X1 U470 ( .A(n392), .B(n530), .ZN(n531) );
  XNOR2_X1 U471 ( .A(n388), .B(n386), .ZN(n385) );
  XNOR2_X1 U472 ( .A(n618), .B(n387), .ZN(n386) );
  XNOR2_X1 U473 ( .A(n390), .B(n389), .ZN(n602) );
  INV_X1 U474 ( .A(KEYINPUT111), .ZN(n389) );
  NAND2_X1 U475 ( .A1(n391), .A2(n415), .ZN(n390) );
  NAND2_X1 U476 ( .A1(n418), .A2(n417), .ZN(n415) );
  NAND2_X1 U477 ( .A1(n567), .A2(n361), .ZN(n563) );
  AND2_X1 U478 ( .A1(n589), .A2(n604), .ZN(n590) );
  INV_X1 U479 ( .A(KEYINPUT60), .ZN(n364) );
  NOR2_X1 U480 ( .A1(n553), .A2(n552), .ZN(n358) );
  INV_X1 U481 ( .A(n650), .ZN(n434) );
  NAND2_X1 U482 ( .A1(n385), .A2(n619), .ZN(n650) );
  NAND2_X1 U483 ( .A1(n689), .A2(n692), .ZN(n359) );
  AND2_X1 U484 ( .A1(n655), .A2(n648), .ZN(n360) );
  AND2_X1 U485 ( .A1(n561), .A2(n698), .ZN(n361) );
  OR2_X1 U486 ( .A1(n575), .A2(G900), .ZN(n362) );
  BUF_X1 U487 ( .A(n546), .Z(n703) );
  XOR2_X1 U488 ( .A(KEYINPUT71), .B(KEYINPUT22), .Z(n363) );
  INV_X1 U489 ( .A(KEYINPUT48), .ZN(n435) );
  INV_X1 U490 ( .A(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U491 ( .A(n365), .B(n364), .ZN(G60) );
  NAND2_X1 U492 ( .A1(n645), .A2(n663), .ZN(n365) );
  NAND2_X1 U493 ( .A1(n366), .A2(n376), .ZN(n383) );
  NOR2_X1 U494 ( .A1(n628), .A2(KEYINPUT2), .ZN(n629) );
  NOR2_X2 U495 ( .A1(n555), .A2(n730), .ZN(n514) );
  XNOR2_X2 U496 ( .A(n513), .B(KEYINPUT0), .ZN(n555) );
  XNOR2_X1 U497 ( .A(n383), .B(n559), .ZN(n571) );
  NAND2_X1 U498 ( .A1(n412), .A2(n367), .ZN(n405) );
  XNOR2_X1 U499 ( .A(n369), .B(n368), .ZN(n758) );
  INV_X1 U500 ( .A(KEYINPUT124), .ZN(n368) );
  NAND2_X1 U501 ( .A1(n703), .A2(n476), .ZN(n706) );
  NAND2_X1 U502 ( .A1(n633), .A2(n501), .ZN(n372) );
  XNOR2_X1 U503 ( .A(n496), .B(n750), .ZN(n633) );
  OR2_X1 U504 ( .A1(n633), .A2(n373), .ZN(n370) );
  NAND2_X1 U505 ( .A1(n501), .A2(n573), .ZN(n375) );
  NAND2_X1 U506 ( .A1(n551), .A2(n359), .ZN(n384) );
  NAND2_X1 U507 ( .A1(n657), .A2(n381), .ZN(n380) );
  AND2_X1 U508 ( .A1(n542), .A2(KEYINPUT44), .ZN(n381) );
  NAND2_X1 U509 ( .A1(n568), .A2(KEYINPUT87), .ZN(n382) );
  INV_X1 U510 ( .A(n602), .ZN(n770) );
  NAND2_X1 U511 ( .A1(n529), .A2(G217), .ZN(n392) );
  NAND2_X1 U512 ( .A1(n505), .A2(G234), .ZN(n394) );
  NAND2_X1 U513 ( .A1(n655), .A2(n395), .ZN(n398) );
  AND2_X1 U514 ( .A1(n568), .A2(n648), .ZN(n395) );
  NAND2_X1 U515 ( .A1(n397), .A2(n396), .ZN(n570) );
  NAND2_X1 U516 ( .A1(n360), .A2(KEYINPUT44), .ZN(n396) );
  NAND2_X1 U517 ( .A1(n398), .A2(n569), .ZN(n397) );
  INV_X1 U518 ( .A(n480), .ZN(n492) );
  NOR2_X1 U519 ( .A1(n555), .A2(n554), .ZN(n401) );
  XNOR2_X2 U520 ( .A(n402), .B(KEYINPUT40), .ZN(n656) );
  NAND2_X1 U521 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U522 ( .A1(n407), .A2(n406), .ZN(n615) );
  XNOR2_X2 U523 ( .A(n587), .B(n586), .ZN(n408) );
  NAND2_X1 U524 ( .A1(n408), .A2(n590), .ZN(n591) );
  INV_X1 U525 ( .A(n742), .ZN(n424) );
  NOR2_X1 U526 ( .A1(n615), .A2(KEYINPUT48), .ZN(n413) );
  XNOR2_X1 U527 ( .A(n414), .B(KEYINPUT5), .ZN(n430) );
  INV_X1 U528 ( .A(n582), .ZN(n418) );
  NAND2_X1 U529 ( .A1(n582), .A2(KEYINPUT36), .ZN(n421) );
  NOR2_X1 U530 ( .A1(n582), .A2(n689), .ZN(n617) );
  NAND2_X1 U531 ( .A1(n742), .A2(n423), .ZN(n733) );
  NAND2_X1 U532 ( .A1(n627), .A2(n424), .ZN(n429) );
  INV_X1 U533 ( .A(KEYINPUT45), .ZN(n425) );
  NAND2_X1 U534 ( .A1(n679), .A2(n691), .ZN(n551) );
  NAND2_X1 U535 ( .A1(n547), .A2(n427), .ZN(n426) );
  XNOR2_X1 U536 ( .A(n545), .B(n428), .ZN(n427) );
  INV_X1 U537 ( .A(KEYINPUT101), .ZN(n428) );
  NAND2_X1 U538 ( .A1(n429), .A2(n436), .ZN(n630) );
  AND2_X1 U539 ( .A1(n429), .A2(n733), .ZN(n736) );
  XNOR2_X2 U540 ( .A(n474), .B(n473), .ZN(n546) );
  XNOR2_X1 U541 ( .A(n430), .B(n432), .ZN(n431) );
  XNOR2_X1 U542 ( .A(n431), .B(n465), .ZN(n470) );
  NAND2_X1 U543 ( .A1(n519), .A2(G210), .ZN(n432) );
  NAND2_X1 U544 ( .A1(n597), .A2(n359), .ZN(n600) );
  INV_X1 U545 ( .A(KEYINPUT87), .ZN(n542) );
  INV_X1 U546 ( .A(KEYINPUT106), .ZN(n580) );
  INV_X1 U547 ( .A(n588), .ZN(n606) );
  XNOR2_X1 U548 ( .A(n591), .B(KEYINPUT109), .ZN(n592) );
  XNOR2_X2 U549 ( .A(G143), .B(G128), .ZN(n487) );
  XNOR2_X2 U550 ( .A(n761), .B(G146), .ZN(n471) );
  XOR2_X1 U551 ( .A(n438), .B(KEYINPUT76), .Z(n440) );
  NAND2_X1 U552 ( .A1(G227), .A2(n505), .ZN(n439) );
  XNOR2_X1 U553 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U554 ( .A(n480), .B(n441), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n471), .B(n442), .ZN(n672) );
  NAND2_X1 U556 ( .A1(n672), .A2(n535), .ZN(n444) );
  XNOR2_X1 U557 ( .A(KEYINPUT68), .B(G469), .ZN(n443) );
  XNOR2_X2 U558 ( .A(n444), .B(n443), .ZN(n543) );
  XNOR2_X1 U559 ( .A(n543), .B(KEYINPUT1), .ZN(n556) );
  XNOR2_X1 U560 ( .A(KEYINPUT97), .B(KEYINPUT24), .ZN(n445) );
  XNOR2_X1 U561 ( .A(n516), .B(n445), .ZN(n447) );
  NAND2_X1 U562 ( .A1(n529), .A2(G221), .ZN(n446) );
  XNOR2_X1 U563 ( .A(n447), .B(n446), .ZN(n455) );
  XNOR2_X1 U564 ( .A(G128), .B(G137), .ZN(n449) );
  XNOR2_X1 U565 ( .A(KEYINPUT23), .B(KEYINPUT98), .ZN(n448) );
  XNOR2_X1 U566 ( .A(n449), .B(n448), .ZN(n453) );
  INV_X1 U567 ( .A(G140), .ZN(n450) );
  XNOR2_X1 U568 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U569 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U570 ( .A(n455), .B(n454), .ZN(n651) );
  XOR2_X1 U571 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n457) );
  XNOR2_X1 U572 ( .A(G902), .B(KEYINPUT15), .ZN(n497) );
  NAND2_X1 U573 ( .A1(n497), .A2(G234), .ZN(n456) );
  XNOR2_X1 U574 ( .A(n457), .B(n456), .ZN(n461) );
  AND2_X1 U575 ( .A1(n461), .A2(G217), .ZN(n458) );
  XNOR2_X1 U576 ( .A(n458), .B(KEYINPUT25), .ZN(n459) );
  XNOR2_X2 U577 ( .A(n460), .B(n459), .ZN(n578) );
  NAND2_X1 U578 ( .A1(n461), .A2(G221), .ZN(n464) );
  INV_X1 U579 ( .A(KEYINPUT100), .ZN(n462) );
  XNOR2_X1 U580 ( .A(n462), .B(KEYINPUT21), .ZN(n463) );
  XNOR2_X1 U581 ( .A(n464), .B(n463), .ZN(n694) );
  XNOR2_X1 U582 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U583 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n468) );
  XNOR2_X1 U584 ( .A(n469), .B(n468), .ZN(n495) );
  XNOR2_X1 U585 ( .A(n470), .B(n495), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n472), .B(n471), .ZN(n659) );
  NOR2_X1 U587 ( .A1(n659), .A2(G902), .ZN(n474) );
  INV_X1 U588 ( .A(G472), .ZN(n473) );
  INV_X1 U589 ( .A(n579), .ZN(n475) );
  NAND2_X1 U590 ( .A1(n476), .A2(n475), .ZN(n479) );
  INV_X1 U591 ( .A(KEYINPUT88), .ZN(n477) );
  XNOR2_X1 U592 ( .A(n477), .B(KEYINPUT33), .ZN(n478) );
  XNOR2_X1 U593 ( .A(n482), .B(n481), .ZN(n486) );
  NAND2_X1 U594 ( .A1(n505), .A2(G224), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n486), .B(n485), .ZN(n490) );
  XOR2_X1 U596 ( .A(n487), .B(n488), .Z(n489) );
  XNOR2_X1 U597 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U598 ( .A(n491), .B(n492), .ZN(n496) );
  XNOR2_X1 U599 ( .A(KEYINPUT16), .B(G122), .ZN(n493) );
  XNOR2_X1 U600 ( .A(n493), .B(KEYINPUT72), .ZN(n494) );
  XNOR2_X1 U601 ( .A(n495), .B(n494), .ZN(n750) );
  INV_X1 U602 ( .A(n497), .ZN(n573) );
  INV_X1 U603 ( .A(G237), .ZN(n498) );
  NAND2_X1 U604 ( .A1(n535), .A2(n498), .ZN(n502) );
  NAND2_X1 U605 ( .A1(n502), .A2(G210), .ZN(n500) );
  INV_X1 U606 ( .A(KEYINPUT92), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U608 ( .A1(n502), .A2(G214), .ZN(n503) );
  XNOR2_X1 U609 ( .A(n503), .B(KEYINPUT93), .ZN(n713) );
  INV_X1 U610 ( .A(n713), .ZN(n610) );
  XNOR2_X1 U611 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n504) );
  XNOR2_X2 U612 ( .A(n583), .B(n504), .ZN(n596) );
  NOR2_X1 U613 ( .A1(G898), .A2(n505), .ZN(n506) );
  XNOR2_X1 U614 ( .A(KEYINPUT95), .B(n506), .ZN(n752) );
  NAND2_X1 U615 ( .A1(G234), .A2(G237), .ZN(n507) );
  XNOR2_X1 U616 ( .A(n507), .B(KEYINPUT94), .ZN(n508) );
  XNOR2_X1 U617 ( .A(KEYINPUT14), .B(n508), .ZN(n509) );
  NAND2_X1 U618 ( .A1(n509), .A2(G902), .ZN(n574) );
  OR2_X1 U619 ( .A1(n752), .A2(n574), .ZN(n510) );
  NAND2_X1 U620 ( .A1(G952), .A2(n509), .ZN(n728) );
  OR2_X1 U621 ( .A1(n728), .A2(G953), .ZN(n576) );
  NAND2_X1 U622 ( .A1(n510), .A2(n576), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n511), .B(KEYINPUT96), .ZN(n512) );
  NAND2_X1 U624 ( .A1(n596), .A2(n512), .ZN(n513) );
  XNOR2_X1 U625 ( .A(n514), .B(KEYINPUT34), .ZN(n538) );
  XNOR2_X1 U626 ( .A(n516), .B(n515), .ZN(n759) );
  XOR2_X1 U627 ( .A(G122), .B(G104), .Z(n518) );
  XNOR2_X1 U628 ( .A(n518), .B(n517), .ZN(n523) );
  XOR2_X1 U629 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n521) );
  NAND2_X1 U630 ( .A1(G214), .A2(n519), .ZN(n520) );
  XNOR2_X1 U631 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n759), .B(n524), .ZN(n642) );
  NAND2_X1 U634 ( .A1(n642), .A2(n535), .ZN(n526) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(G475), .Z(n525) );
  XNOR2_X1 U636 ( .A(n526), .B(n525), .ZN(n550) );
  INV_X1 U637 ( .A(n550), .ZN(n553) );
  XOR2_X1 U638 ( .A(KEYINPUT103), .B(G122), .Z(n528) );
  XNOR2_X1 U639 ( .A(n528), .B(n527), .ZN(n532) );
  XOR2_X1 U640 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U641 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U642 ( .A(n534), .B(n533), .ZN(n666) );
  NAND2_X1 U643 ( .A1(n666), .A2(n535), .ZN(n537) );
  INV_X1 U644 ( .A(G478), .ZN(n536) );
  XNOR2_X1 U645 ( .A(n537), .B(n536), .ZN(n552) );
  NAND2_X1 U646 ( .A1(n538), .A2(n358), .ZN(n541) );
  INV_X1 U647 ( .A(KEYINPUT79), .ZN(n539) );
  XNOR2_X1 U648 ( .A(n539), .B(KEYINPUT35), .ZN(n540) );
  XNOR2_X2 U649 ( .A(n541), .B(n540), .ZN(n657) );
  INV_X1 U650 ( .A(n703), .ZN(n547) );
  OR2_X1 U651 ( .A1(n555), .A2(n706), .ZN(n549) );
  INV_X1 U652 ( .A(KEYINPUT31), .ZN(n548) );
  XNOR2_X1 U653 ( .A(n549), .B(n548), .ZN(n691) );
  OR2_X1 U654 ( .A1(n552), .A2(n550), .ZN(n692) );
  AND2_X1 U655 ( .A1(n553), .A2(n552), .ZN(n715) );
  NAND2_X1 U656 ( .A1(n715), .A2(n694), .ZN(n554) );
  XNOR2_X1 U657 ( .A(n578), .B(KEYINPUT104), .ZN(n695) );
  NAND2_X1 U658 ( .A1(n579), .A2(n695), .ZN(n557) );
  BUF_X1 U659 ( .A(n556), .Z(n698) );
  NOR2_X1 U660 ( .A1(n557), .A2(n698), .ZN(n558) );
  NAND2_X1 U661 ( .A1(n567), .A2(n558), .ZN(n649) );
  INV_X1 U662 ( .A(KEYINPUT86), .ZN(n559) );
  INV_X1 U663 ( .A(n695), .ZN(n560) );
  AND2_X1 U664 ( .A1(n579), .A2(n560), .ZN(n561) );
  XNOR2_X1 U665 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n562) );
  INV_X1 U666 ( .A(n578), .ZN(n564) );
  NAND2_X1 U667 ( .A1(n594), .A2(n564), .ZN(n565) );
  NOR2_X1 U668 ( .A1(n565), .A2(n698), .ZN(n566) );
  NAND2_X1 U669 ( .A1(n567), .A2(n566), .ZN(n648) );
  INV_X1 U670 ( .A(KEYINPUT44), .ZN(n569) );
  NAND2_X1 U671 ( .A1(n571), .A2(n570), .ZN(n572) );
  OR2_X1 U672 ( .A1(n505), .A2(n574), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n362), .A2(n576), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n694), .A2(n605), .ZN(n577) );
  OR2_X1 U675 ( .A1(n578), .A2(n577), .ZN(n593) );
  INV_X1 U676 ( .A(n583), .ZN(n584) );
  INV_X1 U677 ( .A(KEYINPUT108), .ZN(n585) );
  AND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n592), .A2(n358), .ZN(n687) );
  NAND2_X1 U680 ( .A1(n612), .A2(n596), .ZN(n683) );
  INV_X1 U681 ( .A(n683), .ZN(n597) );
  NAND2_X1 U682 ( .A1(n600), .A2(KEYINPUT47), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n687), .A2(n598), .ZN(n599) );
  OR2_X1 U684 ( .A1(n600), .A2(KEYINPUT47), .ZN(n601) );
  XNOR2_X1 U685 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n603) );
  AND2_X1 U686 ( .A1(n712), .A2(n605), .ZN(n607) );
  AND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n608) );
  AND2_X1 U688 ( .A1(n712), .A2(n610), .ZN(n717) );
  NAND2_X1 U689 ( .A1(n717), .A2(n715), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT41), .ZN(n709) );
  NAND2_X1 U691 ( .A1(n612), .A2(n709), .ZN(n614) );
  XNOR2_X1 U692 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n713), .A2(n698), .ZN(n616) );
  INV_X1 U694 ( .A(KEYINPUT107), .ZN(n618) );
  INV_X1 U695 ( .A(n604), .ZN(n619) );
  INV_X1 U696 ( .A(KEYINPUT84), .ZN(n620) );
  OR2_X1 U697 ( .A1(n354), .A2(n692), .ZN(n646) );
  INV_X1 U698 ( .A(KEYINPUT81), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n646), .A2(KEYINPUT2), .ZN(n624) );
  AND2_X1 U700 ( .A1(n624), .A2(KEYINPUT81), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n623), .A2(n625), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n734), .B(KEYINPUT75), .ZN(n628) );
  NOR2_X2 U703 ( .A1(n630), .A2(n629), .ZN(n632) );
  XNOR2_X2 U704 ( .A(n632), .B(n631), .ZN(n658) );
  NAND2_X1 U705 ( .A1(n658), .A2(G210), .ZN(n637) );
  XNOR2_X1 U706 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(KEYINPUT55), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n633), .B(n635), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U710 ( .A(G952), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n638), .A2(G953), .ZN(n663) );
  NAND2_X1 U712 ( .A1(n639), .A2(n663), .ZN(n641) );
  INV_X1 U713 ( .A(KEYINPUT56), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n658), .A2(G475), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n646), .B(G134), .ZN(G36) );
  XNOR2_X1 U718 ( .A(n647), .B(G137), .ZN(G39) );
  XNOR2_X1 U719 ( .A(n648), .B(G110), .ZN(G12) );
  XNOR2_X1 U720 ( .A(n649), .B(G101), .ZN(G3) );
  XNOR2_X1 U721 ( .A(n650), .B(G140), .ZN(G42) );
  BUF_X1 U722 ( .A(n658), .Z(n670) );
  NAND2_X1 U723 ( .A1(n670), .A2(G217), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  INV_X1 U725 ( .A(n663), .ZN(n675) );
  NOR2_X1 U726 ( .A1(n653), .A2(n675), .ZN(G66) );
  XOR2_X1 U727 ( .A(G119), .B(KEYINPUT127), .Z(n654) );
  XNOR2_X1 U728 ( .A(n655), .B(n654), .ZN(G21) );
  XNOR2_X1 U729 ( .A(n656), .B(G131), .ZN(G33) );
  XOR2_X1 U730 ( .A(n657), .B(G122), .Z(G24) );
  NAND2_X1 U731 ( .A1(n658), .A2(G472), .ZN(n662) );
  XOR2_X1 U732 ( .A(KEYINPUT90), .B(KEYINPUT62), .Z(n660) );
  XNOR2_X1 U733 ( .A(n659), .B(n660), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n670), .A2(G478), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT120), .B(n666), .Z(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n669), .A2(n675), .ZN(G63) );
  NAND2_X1 U741 ( .A1(n670), .A2(G469), .ZN(n674) );
  XNOR2_X1 U742 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(G54) );
  NOR2_X1 U746 ( .A1(n357), .A2(n689), .ZN(n677) );
  XOR2_X1 U747 ( .A(KEYINPUT112), .B(n677), .Z(n678) );
  XNOR2_X1 U748 ( .A(G104), .B(n678), .ZN(G6) );
  NOR2_X1 U749 ( .A1(n357), .A2(n692), .ZN(n681) );
  XNOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(G107), .B(n682), .ZN(G9) );
  XOR2_X1 U753 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n685) );
  OR2_X1 U754 ( .A1(n683), .A2(n692), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(n686) );
  XOR2_X1 U756 ( .A(G128), .B(n686), .Z(G30) );
  XNOR2_X1 U757 ( .A(G143), .B(n687), .ZN(G45) );
  OR2_X1 U758 ( .A1(n683), .A2(n689), .ZN(n688) );
  XNOR2_X1 U759 ( .A(G146), .B(n688), .ZN(G48) );
  NOR2_X1 U760 ( .A1(n689), .A2(n691), .ZN(n690) );
  XOR2_X1 U761 ( .A(G113), .B(n690), .Z(G15) );
  NOR2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U763 ( .A(G116), .B(n693), .Z(G18) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U765 ( .A(KEYINPUT49), .B(n696), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U767 ( .A(KEYINPUT114), .B(n699), .Z(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT50), .B(n700), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT115), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U773 ( .A(n708), .B(KEYINPUT51), .ZN(n710) );
  INV_X1 U774 ( .A(n709), .ZN(n729) );
  NOR2_X1 U775 ( .A1(n710), .A2(n729), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n711), .B(KEYINPUT116), .ZN(n725) );
  INV_X1 U777 ( .A(n730), .ZN(n722) );
  INV_X1 U778 ( .A(n712), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U781 ( .A1(n717), .A2(n359), .ZN(n718) );
  XOR2_X1 U782 ( .A(KEYINPUT117), .B(n718), .Z(n719) );
  NAND2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U785 ( .A(KEYINPUT118), .B(n723), .Z(n724) );
  NOR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U787 ( .A(n726), .B(KEYINPUT52), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n734), .A2(n423), .ZN(n735) );
  NAND2_X1 U792 ( .A1(n736), .A2(n735), .ZN(n737) );
  AND2_X1 U793 ( .A1(n737), .A2(n505), .ZN(n738) );
  NAND2_X1 U794 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U795 ( .A(KEYINPUT53), .B(n740), .ZN(n741) );
  XNOR2_X1 U796 ( .A(KEYINPUT119), .B(n741), .ZN(G75) );
  NOR2_X1 U797 ( .A1(n356), .A2(G953), .ZN(n747) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U800 ( .A1(n744), .A2(G898), .ZN(n745) );
  XNOR2_X1 U801 ( .A(n745), .B(KEYINPUT121), .ZN(n746) );
  NOR2_X1 U802 ( .A1(n747), .A2(n746), .ZN(n756) );
  XOR2_X1 U803 ( .A(KEYINPUT122), .B(n748), .Z(n749) );
  XNOR2_X1 U804 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U805 ( .A(G101), .B(n751), .ZN(n753) );
  NAND2_X1 U806 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U807 ( .A(n754), .B(KEYINPUT123), .ZN(n755) );
  XOR2_X1 U808 ( .A(n756), .B(n755), .Z(G69) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n761), .B(n760), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n757), .B(n764), .ZN(n762) );
  NOR2_X1 U812 ( .A1(n762), .A2(G953), .ZN(n763) );
  XNOR2_X1 U813 ( .A(KEYINPUT125), .B(n763), .ZN(n769) );
  XNOR2_X1 U814 ( .A(n764), .B(G227), .ZN(n765) );
  XNOR2_X1 U815 ( .A(n765), .B(KEYINPUT126), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U817 ( .A1(n767), .A2(G953), .ZN(n768) );
  NAND2_X1 U818 ( .A1(n769), .A2(n768), .ZN(G72) );
  XNOR2_X1 U819 ( .A(G125), .B(n770), .ZN(n771) );
  XNOR2_X1 U820 ( .A(n771), .B(KEYINPUT37), .ZN(G27) );
endmodule

