//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT0), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT0), .B(G128), .Z(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n188), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT11), .A2(G134), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G137), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT11), .A2(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT11), .A2(G134), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(G137), .B2(new_n194), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(G137), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n206), .C1(new_n194), .C2(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n203), .A2(new_n208), .A3(KEYINPUT67), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT67), .B1(new_n203), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n193), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n206), .B1(G134), .B2(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n207), .B2(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT65), .B(new_n212), .C1(new_n207), .C2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n190), .A2(new_n218), .A3(G143), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n220), .B(G146), .C1(new_n190), .C2(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n215), .A2(new_n208), .A3(new_n216), .A4(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n211), .A2(KEYINPUT30), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT66), .B(G116), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G119), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT2), .B(G113), .Z(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n196), .A2(new_n198), .ZN(new_n235));
  INV_X1    g049(.A(new_n194), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n206), .B1(new_n237), .B2(new_n205), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n199), .A2(new_n202), .A3(G131), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n193), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n226), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT30), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n227), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n227), .B2(new_n243), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT31), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(G101), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n250), .B(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n211), .A2(new_n226), .A3(new_n234), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n247), .A2(new_n248), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n227), .A2(new_n243), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n227), .A2(new_n243), .A3(new_n244), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n253), .A3(new_n254), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT31), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n241), .A2(new_n233), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  INV_X1    g076(.A(new_n226), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n238), .B2(new_n239), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n203), .A2(new_n208), .A3(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n263), .B1(new_n267), .B2(new_n193), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n262), .B1(new_n268), .B2(new_n234), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n261), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n253), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(KEYINPUT69), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n274));
  INV_X1    g088(.A(new_n261), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n268), .A2(new_n262), .A3(new_n234), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n274), .B1(new_n278), .B2(new_n253), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n255), .A2(new_n260), .A3(new_n273), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NOR2_X1   g095(.A1(G472), .A2(G902), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n254), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n245), .A2(new_n246), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT70), .B1(new_n288), .B2(new_n253), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n257), .A2(new_n254), .A3(new_n258), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n272), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n278), .B2(new_n253), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n268), .A2(new_n234), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n269), .B2(new_n270), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n253), .A2(KEYINPUT29), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(G472), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n187), .B1(new_n286), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT16), .ZN(new_n303));
  XNOR2_X1  g117(.A(G125), .B(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n303), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n303), .A2(new_n306), .A3(G125), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n218), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n304), .B2(KEYINPUT72), .ZN(new_n314));
  OAI211_X1 g128(.A(G146), .B(new_n311), .C1(new_n314), .C2(new_n303), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n317), .A2(new_n190), .A3(G119), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(G119), .B2(new_n190), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n318), .A2(new_n319), .B1(G119), .B2(new_n190), .ZN(new_n320));
  XNOR2_X1  g134(.A(G119), .B(G128), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT24), .B(G110), .Z(new_n322));
  AOI22_X1  g136(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n304), .A2(new_n218), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n315), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(G137), .ZN(new_n331));
  INV_X1    g145(.A(G221), .ZN(new_n332));
  INV_X1    g146(.A(G234), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n332), .A2(new_n333), .A3(G953), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n331), .B(new_n334), .Z(new_n335));
  NAND3_X1  g149(.A1(new_n326), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n324), .A2(new_n325), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT73), .B1(new_n316), .B2(new_n323), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n335), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT25), .B1(new_n342), .B2(G902), .ZN(new_n343));
  INV_X1    g157(.A(G217), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(G234), .B2(new_n295), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n336), .A2(new_n341), .A3(new_n346), .A4(new_n295), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n345), .A2(G902), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n336), .A2(new_n341), .A3(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n255), .A2(new_n260), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n273), .A2(new_n279), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n282), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n283), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n300), .A2(G472), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n302), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G214), .B1(G237), .B2(G902), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT83), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(G110), .B(G122), .Z(new_n367));
  INV_X1    g181(.A(G104), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(new_n368), .B2(G107), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G101), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n369), .A2(new_n372), .A3(new_n376), .A4(new_n373), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n375), .A2(KEYINPUT76), .A3(KEYINPUT4), .A4(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n377), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n375), .B2(KEYINPUT4), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n233), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n371), .A3(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT77), .B1(new_n371), .B2(G104), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n368), .A2(G107), .ZN(new_n388));
  OAI211_X1 g202(.A(G101), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n389), .A2(new_n377), .A3(KEYINPUT78), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT78), .B1(new_n389), .B2(new_n377), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n231), .A2(new_n232), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n228), .A2(KEYINPUT5), .A3(G119), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(G113), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n367), .B1(new_n384), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n367), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n383), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT6), .ZN(new_n402));
  INV_X1    g216(.A(G125), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n193), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n405));
  OR3_X1    g219(.A1(new_n193), .A2(KEYINPUT84), .A3(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(new_n225), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n403), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G224), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G953), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n367), .C1(new_n384), .C2(new_n398), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n402), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n409), .ZN(new_n416));
  INV_X1    g230(.A(new_n411), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT7), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n367), .B(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n396), .A2(new_n393), .B1(new_n377), .B2(new_n389), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n398), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(KEYINPUT7), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n408), .B(KEYINPUT86), .ZN(new_n424));
  INV_X1    g238(.A(new_n404), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n418), .A2(new_n422), .A3(new_n401), .A4(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n415), .A2(new_n295), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT87), .Z(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT88), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n430), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n415), .A2(new_n295), .A3(new_n433), .A4(new_n427), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n366), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(KEYINPUT93), .A2(G952), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT93), .A2(G952), .ZN(new_n437));
  AOI21_X1  g251(.A(G953), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G237), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n333), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G953), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n295), .B(new_n444), .C1(G234), .C2(G237), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G475), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n251), .A2(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n220), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G131), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n206), .A3(new_n451), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(KEYINPUT17), .A3(G131), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n313), .A2(new_n456), .A3(new_n315), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n452), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n314), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n327), .B1(new_n461), .B2(new_n218), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G113), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n368), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT89), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n458), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n458), .A2(new_n463), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(new_n465), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n448), .B1(new_n469), .B2(new_n295), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n453), .A2(new_n455), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n304), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n461), .B2(new_n472), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n315), .B(new_n471), .C1(new_n474), .C2(G146), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n475), .A2(new_n463), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n467), .B1(new_n476), .B2(new_n465), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n448), .A4(new_n295), .ZN(new_n479));
  INV_X1    g293(.A(new_n467), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n465), .B1(new_n475), .B2(new_n463), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n448), .B(new_n295), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT20), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n470), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT9), .B(G234), .Z(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(G217), .A3(new_n444), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n230), .A2(G122), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT90), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n228), .A2(G122), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n230), .A2(new_n490), .A3(G122), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(KEYINPUT14), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(G107), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n220), .A2(G128), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n190), .A2(G143), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT91), .B1(new_n190), .B2(G143), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(G134), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(G107), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n488), .A2(new_n489), .A3(new_n502), .A4(new_n491), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n492), .A2(G107), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n488), .A2(new_n371), .A3(new_n489), .A4(new_n491), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n498), .A2(new_n499), .ZN(new_n507));
  OAI21_X1  g321(.A(G134), .B1(new_n507), .B2(KEYINPUT13), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n500), .ZN(new_n509));
  INV_X1    g323(.A(new_n507), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT13), .A3(G134), .A4(new_n495), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n505), .A2(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n486), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n514));
  INV_X1    g328(.A(new_n486), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n505), .A2(new_n506), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n509), .A2(new_n511), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G478), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n519), .A2(new_n520), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n521), .B1(new_n525), .B2(new_n523), .ZN(new_n526));
  AND4_X1   g340(.A1(new_n447), .A2(new_n484), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n435), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n332), .B1(new_n485), .B2(new_n295), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G140), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n444), .A2(G227), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n392), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n225), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n389), .A2(new_n377), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT78), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n389), .A2(new_n377), .A3(KEYINPUT78), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT79), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n407), .A2(new_n537), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT10), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n382), .B2(new_n193), .ZN(new_n547));
  INV_X1    g361(.A(new_n267), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n544), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n535), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n534), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT80), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT12), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n225), .B1(new_n539), .B2(new_n540), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(new_n545), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n238), .A2(new_n239), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT12), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n545), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(KEYINPUT80), .C1(new_n392), .C2(new_n225), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n564), .A3(new_n267), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT82), .B(new_n535), .C1(new_n549), .C2(new_n550), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n553), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n295), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT81), .B1(new_n566), .B2(new_n549), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT81), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n554), .A2(new_n562), .A3(new_n573), .A4(new_n565), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n574), .A3(new_n535), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n555), .A2(new_n550), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(G469), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(G469), .A2(G902), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n528), .A2(new_n529), .A3(new_n531), .A4(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n579), .A2(new_n435), .A3(new_n531), .A4(new_n527), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT94), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n363), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(new_n376), .ZN(G3));
  AND2_X1   g399(.A1(new_n579), .A2(new_n531), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n280), .A2(new_n295), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G472), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(new_n358), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n589), .A3(new_n355), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n513), .A2(new_n518), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT33), .Z(new_n592));
  OAI21_X1  g406(.A(G478), .B1(new_n592), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n484), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n519), .A2(new_n522), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n364), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n428), .A2(new_n430), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(new_n434), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n447), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT34), .B(G104), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  INV_X1    g418(.A(new_n470), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n479), .A2(new_n483), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n524), .A2(new_n526), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n446), .B(KEYINPUT96), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n600), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n590), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT35), .B(G107), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  NOR2_X1   g428(.A1(new_n340), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n339), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n351), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n348), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n588), .A2(new_n618), .A3(new_n358), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n588), .A2(new_n618), .A3(KEYINPUT97), .A4(new_n358), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n580), .A2(new_n582), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT37), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G110), .ZN(G12));
  AND3_X1   g439(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n361), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT71), .B1(new_n360), .B2(new_n361), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n441), .B1(new_n629), .B2(new_n445), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n609), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n631), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n632), .A2(new_n600), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n628), .A2(new_n586), .A3(new_n618), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  XOR2_X1   g452(.A(new_n630), .B(KEYINPUT39), .Z(new_n639));
  NAND2_X1  g453(.A1(new_n586), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT40), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n618), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n287), .A2(new_n253), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n646), .B2(new_n296), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n288), .B2(new_n272), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G472), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n360), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n360), .A2(KEYINPUT99), .A3(new_n649), .ZN(new_n653));
  INV_X1    g467(.A(new_n608), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n484), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n432), .A2(new_n434), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n645), .A2(new_n656), .A3(new_n364), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NAND2_X1  g474(.A1(G478), .A2(G902), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n591), .B(KEYINPUT33), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n595), .B(new_n661), .C1(new_n662), .C2(new_n522), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n663), .A2(new_n484), .A3(new_n630), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n600), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT100), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n628), .A2(new_n586), .A3(new_n618), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G146), .ZN(G48));
  NOR3_X1   g482(.A1(new_n626), .A2(new_n627), .A3(new_n354), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  INV_X1    g484(.A(new_n601), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n569), .A2(new_n295), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G469), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(KEYINPUT101), .A3(new_n571), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n675), .A3(G469), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n530), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n302), .A2(new_n677), .A3(new_n355), .A4(new_n362), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT102), .B1(new_n679), .B2(new_n601), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT41), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G113), .ZN(G15));
  NOR2_X1   g497(.A1(new_n679), .A2(new_n611), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n228), .ZN(G18));
  AND4_X1   g499(.A1(new_n302), .A2(new_n362), .A3(new_n527), .A4(new_n618), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n677), .A2(new_n600), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  AOI22_X1  g503(.A1(new_n259), .A2(KEYINPUT31), .B1(new_n297), .B2(new_n272), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n255), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n282), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n355), .A2(new_n588), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT104), .Z(new_n696));
  AND2_X1   g510(.A1(new_n655), .A2(new_n610), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n687), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  INV_X1    g513(.A(new_n664), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n694), .A2(new_n588), .A3(new_n618), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT105), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n694), .A2(new_n588), .A3(new_n703), .A4(new_n618), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n687), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NAND2_X1  g521(.A1(new_n577), .A2(KEYINPUT106), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n575), .A2(new_n709), .A3(G469), .A4(new_n576), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n571), .A3(new_n578), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n657), .A2(new_n598), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n531), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n664), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n302), .A2(new_n713), .A3(new_n355), .A4(new_n362), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(new_n700), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(KEYINPUT107), .B(new_n718), .C1(new_n719), .C2(new_n700), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n717), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n726), .B(new_n717), .C1(new_n722), .C2(new_n723), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND4_X1  g544(.A1(new_n669), .A2(new_n635), .A3(new_n632), .A4(new_n713), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n575), .A2(new_n576), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n733), .B(G469), .C1(new_n734), .C2(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g550(.A1(KEYINPUT45), .A2(G469), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n577), .A2(KEYINPUT109), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n578), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n578), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n571), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n531), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n639), .ZN(new_n747));
  INV_X1    g561(.A(new_n712), .ZN(new_n748));
  INV_X1    g562(.A(new_n589), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n663), .A2(new_n594), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n757), .A3(new_n618), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n748), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n747), .B(new_n760), .C1(new_n759), .C2(new_n758), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  NAND2_X1  g576(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n745), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n700), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n628), .A2(new_n748), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n354), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  AND2_X1   g583(.A1(new_n696), .A2(new_n687), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n440), .B1(new_n754), .B2(new_n756), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n674), .A2(new_n676), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n530), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n765), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n696), .A3(new_n712), .A4(new_n771), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n354), .B1(new_n652), .B2(new_n653), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n531), .A2(new_n773), .A3(new_n441), .A4(new_n712), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT119), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n484), .A3(new_n663), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n677), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n658), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n696), .A2(new_n787), .A3(new_n771), .A4(new_n598), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(KEYINPUT50), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(KEYINPUT50), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n778), .A2(new_n757), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n702), .A2(new_n704), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n783), .A2(new_n784), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n776), .A2(new_n785), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT51), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n438), .B(new_n772), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n780), .A2(new_n597), .A3(new_n782), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n770), .A2(new_n697), .B1(new_n678), .B2(new_n680), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n608), .A2(new_n484), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n596), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n805), .A2(new_n435), .A3(new_n610), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n586), .A3(new_n589), .A4(new_n355), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n623), .B(new_n807), .C1(new_n363), .C2(new_n583), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n792), .B2(new_n714), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n302), .A2(new_n362), .A3(new_n586), .A4(new_n618), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n654), .A2(new_n607), .A3(new_n606), .A4(new_n631), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT112), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n748), .B1(new_n811), .B2(KEYINPUT112), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(new_n731), .ZN(new_n815));
  INV_X1    g629(.A(new_n611), .ZN(new_n816));
  INV_X1    g630(.A(new_n679), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n816), .A2(new_n817), .B1(new_n686), .B2(new_n687), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n803), .A2(new_n809), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n725), .B2(new_n728), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n618), .B1(new_n822), .B2(new_n630), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n631), .A2(KEYINPUT113), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n823), .A2(new_n711), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n655), .A2(new_n600), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n531), .A3(new_n650), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n637), .A2(new_n667), .A3(new_n706), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n810), .A2(new_n636), .B1(new_n687), .B2(new_n705), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n667), .A4(new_n827), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n828), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT114), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n828), .A2(new_n837), .A3(new_n830), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n820), .A2(new_n821), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n830), .B1(new_n829), .B2(new_n833), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n681), .A2(new_n818), .A3(new_n698), .ZN(new_n844));
  INV_X1    g658(.A(new_n808), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n714), .A2(new_n792), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n731), .A3(new_n846), .A4(new_n814), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n727), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT53), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n840), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n821), .B1(new_n843), .B2(new_n850), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n844), .B(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n724), .A2(new_n847), .A3(new_n821), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n839), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n852), .A2(new_n859), .A3(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n791), .A2(new_n715), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT48), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n802), .A2(new_n862), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(G952), .A2(G953), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n773), .B(KEYINPUT49), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n658), .A2(new_n530), .A3(new_n366), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n777), .A2(new_n869), .A3(new_n750), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT111), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(G75));
  AOI21_X1  g687(.A(new_n295), .B1(new_n853), .B2(new_n858), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT56), .B1(new_n874), .B2(new_n430), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n402), .A2(new_n414), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(new_n412), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT55), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(KEYINPUT121), .ZN(new_n880));
  AOI211_X1 g694(.A(KEYINPUT56), .B(new_n880), .C1(new_n874), .C2(new_n431), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n444), .A2(G952), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(G51));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n739), .B(KEYINPUT122), .Z(new_n885));
  AOI211_X1 g699(.A(new_n295), .B(new_n885), .C1(new_n853), .C2(new_n858), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n578), .B(KEYINPUT57), .Z(new_n887));
  AND3_X1   g701(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n854), .B1(new_n853), .B2(new_n858), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n886), .B1(new_n890), .B2(new_n569), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n884), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  INV_X1    g706(.A(new_n882), .ZN(new_n893));
  INV_X1    g707(.A(new_n569), .ZN(new_n894));
  INV_X1    g708(.A(new_n842), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n834), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n820), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n839), .A2(new_n856), .A3(new_n857), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n859), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n894), .B1(new_n900), .B2(new_n887), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT123), .B(new_n893), .C1(new_n901), .C2(new_n886), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n892), .A2(new_n902), .ZN(G54));
  NAND3_X1  g717(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n904));
  INV_X1    g718(.A(new_n477), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n882), .ZN(G60));
  XOR2_X1   g722(.A(new_n661), .B(KEYINPUT59), .Z(new_n909));
  AOI211_X1 g723(.A(new_n592), .B(new_n909), .C1(new_n899), .C2(new_n859), .ZN(new_n910));
  INV_X1    g724(.A(new_n909), .ZN(new_n911));
  INV_X1    g725(.A(new_n863), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT117), .B1(new_n852), .B2(new_n859), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n882), .B(new_n910), .C1(new_n914), .C2(new_n592), .ZN(G63));
  NAND2_X1  g729(.A1(new_n853), .A2(new_n858), .ZN(new_n916));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n350), .A2(new_n352), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n616), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n921), .B(new_n893), .C1(new_n922), .C2(new_n919), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n443), .B2(new_n410), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n844), .A2(new_n808), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n876), .B1(G898), .B2(new_n444), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G69));
  NAND3_X1  g745(.A1(new_n747), .A2(new_n715), .A3(new_n826), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n731), .A2(new_n768), .A3(new_n761), .A4(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n831), .A2(new_n667), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n729), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n444), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n241), .A2(new_n242), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n227), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n474), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n629), .B2(G953), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n444), .B1(G227), .B2(G900), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT127), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n944), .A2(KEYINPUT127), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n934), .A2(new_n659), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n669), .A2(new_n641), .A3(new_n712), .A4(new_n805), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT125), .Z(new_n950));
  NAND3_X1  g764(.A1(new_n768), .A2(new_n761), .A3(new_n950), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT126), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(new_n948), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n444), .A3(new_n940), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n943), .A2(new_n945), .A3(new_n946), .A4(new_n955), .ZN(new_n956));
  AOI211_X1 g770(.A(G953), .B(new_n939), .C1(new_n952), .C2(new_n953), .ZN(new_n957));
  OAI211_X1 g771(.A(KEYINPUT127), .B(new_n944), .C1(new_n957), .C2(new_n942), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(G72));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  INV_X1    g775(.A(new_n927), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n954), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n253), .A3(new_n290), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n935), .B2(new_n962), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n272), .A3(new_n288), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n289), .A2(new_n259), .A3(new_n292), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n840), .A2(new_n851), .A3(new_n961), .A4(new_n967), .ZN(new_n968));
  AND4_X1   g782(.A1(new_n893), .A2(new_n964), .A3(new_n966), .A4(new_n968), .ZN(G57));
endmodule


