//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n203), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n203), .A2(new_n207), .B1(KEYINPUT16), .B2(new_n204), .ZN(new_n209));
  OAI21_X1  g008(.A(G8gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n203), .A2(new_n204), .A3(new_n207), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n203), .A2(new_n207), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G43gat), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(G43gat), .A2(G50gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT88), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n219), .A2(KEYINPUT88), .A3(new_n220), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227));
  INV_X1    g026(.A(G36gat), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G29gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n219), .A2(new_n221), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n231), .A2(new_n233), .B1(new_n234), .B2(KEYINPUT15), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n234), .A3(KEYINPUT15), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n227), .B1(new_n226), .B2(new_n235), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT17), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n237), .A4(new_n236), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n216), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n238), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n247), .A2(new_n241), .B1(new_n210), .B2(new_n215), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n244), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT91), .B1(new_n249), .B2(KEYINPUT18), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n240), .A2(new_n243), .ZN(new_n251));
  INV_X1    g050(.A(new_n216), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n248), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n245), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n253), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n254), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n245), .B(KEYINPUT13), .Z(new_n261));
  NOR3_X1   g060(.A1(new_n216), .A2(new_n239), .A3(new_n238), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n248), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G141gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G197gat), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT11), .B(G169gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n257), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n263), .A3(new_n260), .ZN(new_n272));
  INV_X1    g071(.A(new_n268), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n259), .A2(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G228gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G141gat), .B(G148gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT2), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n280), .A2(KEYINPUT74), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(KEYINPUT74), .B2(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  OR2_X1    g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n280), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n288), .B2(KEYINPUT2), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n280), .A2(new_n290), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n279), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(KEYINPUT22), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n294), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n289), .A2(KEYINPUT77), .A3(new_n294), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n296), .B1(new_n304), .B2(new_n279), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n277), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n277), .B1(new_n297), .B2(new_n305), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n304), .A2(KEYINPUT29), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n316), .A2(KEYINPUT81), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT3), .B1(new_n316), .B2(KEYINPUT81), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n295), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OR3_X1    g118(.A1(new_n315), .A2(KEYINPUT82), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT82), .B1(new_n315), .B2(new_n319), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G22gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n323), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(new_n218), .ZN(new_n329));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  NAND4_X1  g130(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n326), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n327), .B1(new_n322), .B2(new_n323), .ZN(new_n334));
  INV_X1    g133(.A(new_n331), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n333), .A2(new_n324), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n295), .A2(new_n296), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT1), .ZN(new_n341));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  INV_X1    g146(.A(new_n343), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n307), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n309), .A2(KEYINPUT4), .A3(new_n343), .A4(new_n310), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n338), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n346), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n339), .B2(new_n344), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(KEYINPUT78), .A3(new_n351), .A4(new_n349), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n307), .B(new_n348), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n354), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT0), .ZN(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  NAND4_X1  g164(.A1(new_n309), .A2(new_n347), .A3(new_n343), .A4(new_n310), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT4), .B1(new_n307), .B2(new_n348), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(new_n358), .A3(new_n355), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n361), .A2(new_n369), .ZN(new_n371));
  INV_X1    g170(.A(new_n365), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT6), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(new_n372), .ZN(new_n374));
  INV_X1    g173(.A(new_n360), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n353), .B2(new_n356), .ZN(new_n376));
  INV_X1    g175(.A(new_n369), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT6), .B(new_n372), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n370), .A2(new_n373), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G169gat), .ZN(new_n384));
  INV_X1    g183(.A(G176gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n386), .A2(KEYINPUT26), .A3(new_n387), .ZN(new_n388));
  AOI211_X1 g187(.A(new_n383), .B(new_n388), .C1(KEYINPUT26), .C2(new_n387), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT27), .B(G183gat), .ZN(new_n390));
  INV_X1    g189(.A(G190gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT28), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n383), .A2(KEYINPUT24), .ZN(new_n397));
  NAND2_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n398));
  MUX2_X1   g197(.A(G183gat), .B(new_n398), .S(G190gat), .Z(new_n399));
  AND2_X1   g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n387), .A2(KEYINPUT23), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT23), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n401), .B(new_n403), .C1(new_n384), .C2(new_n385), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n396), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n396), .ZN(new_n406));
  AND2_X1   g205(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n382), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n399), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n413), .B(KEYINPUT72), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n395), .B2(new_n411), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n415), .B(new_n305), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n412), .B2(new_n278), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n412), .B2(new_n414), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n419), .B2(new_n305), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n424), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n427));
  OR3_X1    g226(.A1(new_n420), .A2(KEYINPUT30), .A3(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n337), .B1(new_n381), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n348), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n395), .A2(new_n411), .A3(new_n343), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n432), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n437), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT66), .B(new_n439), .C1(new_n433), .C2(new_n434), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT32), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(new_n438), .B2(new_n440), .ZN(new_n443));
  XNOR2_X1  g242(.A(G15gat), .B(G43gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT67), .ZN(new_n445));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n441), .A2(new_n443), .A3(KEYINPUT68), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n441), .B1(KEYINPUT33), .B2(new_n447), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n435), .A2(KEYINPUT34), .A3(new_n437), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT70), .ZN(new_n458));
  INV_X1    g257(.A(new_n435), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n436), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(KEYINPUT70), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n456), .B1(new_n463), .B2(KEYINPUT71), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n453), .B1(new_n450), .B2(new_n451), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT71), .B1(new_n466), .B2(new_n456), .ZN(new_n467));
  INV_X1    g266(.A(new_n463), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n465), .B(KEYINPUT36), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n468), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n466), .A2(new_n463), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n431), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n431), .A2(new_n476), .A3(new_n473), .A4(new_n469), .ZN(new_n477));
  INV_X1    g276(.A(new_n337), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n368), .A2(new_n345), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n354), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n365), .B1(new_n480), .B2(KEYINPUT39), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT39), .B1(new_n359), .B2(new_n354), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT85), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(KEYINPUT40), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n484), .B(new_n486), .Z(new_n487));
  NAND2_X1  g286(.A1(new_n371), .A2(new_n372), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n430), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n373), .A2(new_n370), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n374), .A2(new_n380), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n424), .B1(new_n420), .B2(KEYINPUT37), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n415), .B(new_n304), .C1(new_n414), .C2(new_n416), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(KEYINPUT37), .C1(new_n419), .C2(new_n304), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(KEYINPUT37), .B2(new_n420), .ZN(new_n498));
  OAI221_X1 g297(.A(new_n425), .B1(new_n493), .B2(new_n497), .C1(new_n498), .C2(new_n496), .ZN(new_n499));
  OAI221_X1 g298(.A(new_n478), .B1(new_n487), .B2(new_n489), .C1(new_n492), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n477), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n478), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n492), .A2(new_n429), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT35), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n471), .A2(new_n472), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT87), .B1(new_n381), .B2(new_n430), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n509), .A3(new_n429), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n337), .A2(KEYINPUT35), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n507), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n274), .B1(new_n501), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(G57gat), .A2(G64gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(G57gat), .A2(G64gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518));
  NAND2_X1  g317(.A1(G71gat), .A2(G78gat), .ZN(new_n519));
  INV_X1    g318(.A(G71gat), .ZN(new_n520));
  INV_X1    g319(.A(G78gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT9), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(KEYINPUT93), .A3(new_n516), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n516), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n216), .B1(KEYINPUT21), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G155gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G127gat), .ZN(new_n543));
  XOR2_X1   g342(.A(G183gat), .B(G211gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n538), .A2(new_n545), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n556));
  AND4_X1   g355(.A1(new_n551), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  AND2_X1   g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G99gat), .ZN(new_n562));
  INV_X1    g361(.A(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(KEYINPUT97), .A3(new_n550), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n557), .A2(new_n566), .A3(KEYINPUT98), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT98), .B1(new_n557), .B2(new_n566), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n549), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n561), .A2(new_n565), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n551), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n566), .A3(KEYINPUT98), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT99), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n572), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n251), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n238), .A2(new_n239), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584));
  NOR3_X1   g383(.A1(new_n578), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT96), .Z(new_n588));
  XOR2_X1   g387(.A(G134gat), .B(G162gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n584), .B1(new_n578), .B2(new_n583), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n586), .A2(KEYINPUT100), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n590), .B(KEYINPUT100), .Z(new_n593));
  INV_X1    g392(.A(new_n591), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n594), .B2(new_n585), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n548), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G230gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n276), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n569), .A2(new_n575), .A3(new_n531), .A4(new_n576), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n567), .A2(new_n568), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n571), .A2(new_n604), .A3(new_n572), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT101), .B1(new_n557), .B2(new_n566), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n532), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT10), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n525), .B(KEYINPUT10), .C1(new_n529), .C2(new_n530), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(new_n569), .A3(new_n575), .A4(new_n576), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n601), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n602), .A2(new_n608), .A3(new_n600), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n598), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n492), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n381), .A2(KEYINPUT102), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n514), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g432(.A1(new_n514), .A2(new_n626), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n429), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n211), .B2(new_n635), .ZN(new_n638));
  MUX2_X1   g437(.A(new_n637), .B(new_n638), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g438(.A1(new_n469), .A2(new_n473), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(G15gat), .B1(new_n634), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n506), .A2(G15gat), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n634), .B2(new_n643), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n634), .A2(new_n478), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  NAND2_X1  g446(.A1(new_n501), .A2(new_n513), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n596), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n431), .A2(new_n469), .A3(new_n473), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n505), .A2(new_n512), .B1(new_n652), .B2(new_n500), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(new_n596), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n548), .B(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n656), .A2(new_n274), .A3(new_n623), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n232), .B1(new_n658), .B2(new_n631), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  INV_X1    g460(.A(new_n548), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(new_n596), .A3(new_n623), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n630), .A2(G29gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n514), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n514), .A2(new_n663), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(KEYINPUT45), .A3(new_n664), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n660), .A2(new_n661), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n667), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT104), .B1(new_n671), .B2(new_n659), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(G1328gat));
  AOI21_X1  g472(.A(new_n228), .B1(new_n658), .B2(new_n430), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n514), .A2(new_n228), .A3(new_n430), .A4(new_n663), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT46), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(KEYINPUT46), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n675), .A2(new_n676), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n678), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(new_n681), .B2(new_n674), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n658), .A2(G43gat), .A3(new_n640), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n514), .A2(new_n507), .A3(new_n663), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(new_n217), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1330gat));
  NOR2_X1   g488(.A1(new_n478), .A2(G50gat), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n668), .A2(new_n690), .B1(KEYINPUT107), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n651), .A2(new_n654), .A3(new_n337), .A4(new_n657), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G50gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n691), .A2(KEYINPUT107), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n652), .A2(new_n500), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n513), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n260), .A2(new_n263), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n244), .A2(new_n248), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT18), .B1(new_n701), .B2(new_n245), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n273), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n250), .A2(new_n258), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n269), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n548), .A2(new_n705), .A3(new_n597), .A4(new_n624), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n699), .A2(KEYINPUT108), .A3(new_n706), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n631), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n429), .B(KEYINPUT109), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n717));
  INV_X1    g516(.A(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT110), .Z(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n711), .A2(new_n714), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n709), .A2(new_n710), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT111), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n722), .A2(new_n717), .A3(new_n724), .A4(new_n718), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1333gat));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n520), .A3(new_n507), .ZN(new_n729));
  OAI21_X1  g528(.A(G71gat), .B1(new_n723), .B2(new_n641), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n729), .B2(new_n730), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1334gat));
  NOR2_X1   g533(.A1(new_n723), .A2(new_n478), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n521), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n662), .A2(new_n705), .A3(new_n624), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n651), .A2(new_n654), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738), .B2(new_n630), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n662), .A2(new_n705), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n699), .A2(new_n597), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n597), .A4(new_n740), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n624), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n630), .A2(G85gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(G1336gat));
  NOR2_X1   g547(.A1(new_n715), .A2(G92gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n745), .A2(KEYINPUT113), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G92gat), .B1(new_n738), .B2(new_n715), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(KEYINPUT52), .B(G92gat), .C1(new_n738), .C2(new_n429), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n745), .A2(new_n749), .B1(KEYINPUT113), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n738), .B2(new_n641), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n507), .A2(new_n562), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n746), .B2(new_n758), .ZN(G1338gat));
  NAND4_X1  g558(.A1(new_n651), .A2(new_n654), .A3(new_n337), .A4(new_n737), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n337), .A2(new_n563), .A3(new_n623), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT115), .Z(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n743), .B2(new_n744), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n761), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n760), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n760), .B2(G106gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(new_n764), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n625), .A2(new_n705), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n602), .A2(new_n608), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT10), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n600), .B1(new_n777), .B2(new_n612), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n612), .A2(new_n600), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT54), .B1(new_n609), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n782), .B(new_n601), .C1(new_n609), .C2(new_n613), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n620), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n774), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n779), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n614), .A3(KEYINPUT54), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n620), .A4(new_n783), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(new_n622), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n270), .A2(new_n250), .A3(new_n258), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n262), .A2(new_n248), .ZN(new_n793));
  OAI22_X1  g592(.A1(new_n793), .A2(new_n261), .B1(new_n701), .B2(new_n245), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n267), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n796), .A3(new_n597), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n623), .A3(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n274), .B2(new_n790), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n597), .B1(new_n800), .B2(KEYINPUT117), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n802), .C1(new_n274), .C2(new_n790), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n798), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n655), .B1(new_n804), .B2(KEYINPUT118), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n806), .B(new_n798), .C1(new_n801), .C2(new_n803), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n773), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(new_n337), .A3(new_n630), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n507), .A3(new_n715), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n274), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n502), .A3(new_n715), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n274), .A2(G113gat), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT119), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(G1340gat));
  INV_X1    g615(.A(G120gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n811), .A2(new_n817), .A3(new_n624), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n813), .A2(new_n624), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n817), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n811), .B2(new_n655), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n548), .A2(G127gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n813), .B2(new_n822), .ZN(G1342gat));
  NAND2_X1  g622(.A1(new_n810), .A2(new_n502), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n430), .A2(G134gat), .A3(new_n596), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n824), .A2(KEYINPUT56), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n811), .B2(new_n596), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT56), .B1(new_n824), .B2(new_n825), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G1343gat));
  NAND4_X1  g628(.A1(new_n473), .A2(new_n469), .A3(new_n628), .A4(new_n629), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n809), .A2(new_n478), .A3(new_n716), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n274), .A2(G141gat), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(KEYINPUT58), .ZN(new_n834));
  OR3_X1    g633(.A1(new_n830), .A2(KEYINPUT120), .A3(new_n716), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT120), .B1(new_n830), .B2(new_n716), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(new_n808), .B2(new_n337), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n337), .A2(KEYINPUT57), .ZN(new_n839));
  INV_X1    g638(.A(new_n622), .ZN(new_n840));
  INV_X1    g639(.A(new_n780), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n774), .B1(new_n841), .B2(new_n614), .ZN(new_n842));
  INV_X1    g641(.A(new_n784), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n781), .B2(new_n784), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n705), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n799), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT122), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n850), .A3(new_n799), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n597), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n797), .B1(new_n852), .B2(KEYINPUT123), .ZN(new_n853));
  INV_X1    g652(.A(new_n851), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n847), .B2(new_n799), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT123), .B(new_n596), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n548), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n839), .B1(new_n858), .B2(new_n773), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n837), .B1(new_n838), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G141gat), .B1(new_n860), .B2(new_n274), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n834), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n837), .B(KEYINPUT124), .C1(new_n838), .C2(new_n859), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n705), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n833), .B1(new_n866), .B2(G141gat), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(G1344gat));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(G148gat), .C1(new_n831), .C2(new_n623), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n864), .A2(new_n870), .A3(new_n623), .A4(new_n865), .ZN(new_n872));
  INV_X1    g671(.A(G148gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n809), .A2(new_n839), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n852), .A2(new_n798), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n773), .B1(new_n662), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n337), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n623), .B(new_n837), .C1(new_n874), .C2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n873), .B1(new_n878), .B2(KEYINPUT59), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n871), .B1(new_n872), .B2(new_n879), .ZN(G1345gat));
  INV_X1    g679(.A(G155gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n831), .A2(new_n881), .A3(new_n662), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n864), .A2(new_n656), .A3(new_n865), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n881), .ZN(G1346gat));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n597), .A3(new_n865), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G162gat), .ZN(new_n886));
  INV_X1    g685(.A(new_n830), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n430), .A2(G162gat), .A3(new_n596), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n808), .A2(new_n337), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n809), .A2(new_n337), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n631), .A2(new_n429), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n507), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(new_n384), .A3(new_n274), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n809), .A2(new_n631), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n716), .A2(new_n502), .A3(new_n478), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n705), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n900), .B1(new_n384), .B2(new_n906), .ZN(G1348gat));
  OAI21_X1  g706(.A(G176gat), .B1(new_n899), .B2(new_n624), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n623), .A2(new_n385), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n904), .B2(new_n909), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n899), .B2(new_n655), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n662), .A2(new_n390), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n904), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n905), .A2(new_n391), .A3(new_n597), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n895), .A2(new_n597), .A3(new_n898), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(G190gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n916), .B2(G190gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  INV_X1    g719(.A(new_n896), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n640), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n874), .B2(new_n877), .ZN(new_n923));
  INV_X1    g722(.A(G197gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(new_n274), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n640), .A2(new_n478), .A3(new_n715), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n808), .A2(new_n926), .A3(new_n630), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n705), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n925), .B1(new_n924), .B2(new_n931), .ZN(G1352gat));
  OAI21_X1  g731(.A(G204gat), .B1(new_n923), .B2(new_n624), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n624), .A2(G204gat), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT62), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n927), .A2(KEYINPUT62), .A3(new_n934), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(G1353gat));
  NAND4_X1  g736(.A1(new_n929), .A2(new_n299), .A3(new_n662), .A4(new_n930), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n923), .A2(new_n548), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n923), .B2(new_n596), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n929), .A2(new_n300), .A3(new_n597), .A4(new_n930), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT127), .Z(G1355gat));
endmodule


