//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AND2_X1   g0010(.A1(G77), .A2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G116), .C2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n223), .A2(new_n207), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n225), .B(new_n226), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(G58), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n216), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n219), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n221), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n222), .A2(G1698), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G226), .B2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G97), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n256), .A2(new_n261), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n264), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n252), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n214), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(KEYINPUT13), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n271), .A2(KEYINPUT14), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n270), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(new_n274), .B2(G169), .ZN(new_n278));
  OR3_X1    g0078(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n228), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT69), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n259), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n286), .A2(new_n204), .B1(new_n229), .B2(G68), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n281), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(new_n288), .B(KEYINPUT11), .Z(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G20), .A3(new_n213), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT12), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n280), .B(new_n228), .C1(G1), .C2(new_n229), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n213), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n279), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n271), .A2(G190), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n274), .A2(G200), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT70), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT18), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n257), .B2(G33), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n259), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(G223), .A2(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n220), .A2(G1698), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n264), .ZN(new_n314));
  INV_X1    g0114(.A(new_n254), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n267), .B2(new_n222), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n317), .A3(G179), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n266), .B1(new_n311), .B2(new_n312), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n319), .B2(new_n316), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n259), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT71), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n258), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(new_n229), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT7), .B1(new_n308), .B2(G20), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(G68), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n221), .A2(new_n213), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n231), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n282), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT3), .B(G33), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n324), .B1(new_n335), .B2(G20), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n213), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n334), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n281), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT67), .A2(G58), .ZN(new_n342));
  XOR2_X1   g0142(.A(new_n342), .B(KEYINPUT8), .Z(new_n343));
  MUX2_X1   g0143(.A(new_n294), .B(new_n341), .S(new_n343), .Z(new_n344));
  AOI221_X4 g0144(.A(new_n303), .B1(new_n318), .B2(new_n320), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n340), .A2(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n318), .A2(new_n320), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT18), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(G200), .B1(new_n319), .B2(new_n316), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n314), .A2(new_n317), .A3(G190), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n340), .A2(new_n351), .A3(new_n352), .A4(new_n344), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT17), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n335), .A2(G232), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n335), .A2(G238), .A3(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(new_n215), .C2(new_n335), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n254), .B1(new_n359), .B2(new_n264), .ZN(new_n360));
  INV_X1    g0160(.A(new_n267), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G244), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n275), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT8), .B(G58), .Z(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n286), .ZN(new_n369));
  INV_X1    g0169(.A(new_n341), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n369), .A2(new_n281), .B1(new_n204), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n204), .B2(new_n294), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n365), .B(new_n372), .C1(G169), .C2(new_n364), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n355), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n376));
  OAI211_X1 g0176(.A(KEYINPUT70), .B(new_n301), .C1(new_n376), .C2(new_n296), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n335), .A2(G222), .A3(new_n356), .ZN(new_n379));
  XOR2_X1   g0179(.A(new_n379), .B(KEYINPUT66), .Z(new_n380));
  NAND3_X1  g0180(.A1(new_n335), .A2(G223), .A3(G1698), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n204), .B2(new_n335), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n264), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n361), .A2(G226), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n315), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G190), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n203), .A2(new_n229), .ZN(new_n387));
  INV_X1    g0187(.A(G150), .ZN(new_n388));
  INV_X1    g0188(.A(new_n282), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n343), .A2(new_n286), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n281), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n294), .A2(new_n219), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n370), .A2(new_n219), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT9), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n383), .A2(new_n384), .A3(new_n315), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n386), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT10), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n385), .A2(new_n275), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(new_n394), .C1(G169), .C2(new_n385), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n364), .A2(KEYINPUT68), .A3(G190), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT68), .ZN(new_n403));
  INV_X1    g0203(.A(G190), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n363), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n372), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n363), .A2(G200), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n399), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  OR3_X1    g0209(.A1(new_n302), .A2(new_n378), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(G244), .B(new_n258), .C1(new_n321), .C2(new_n322), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT4), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n258), .A2(new_n260), .A3(G250), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT4), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G283), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n335), .A2(KEYINPUT4), .A3(G244), .A4(new_n356), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n413), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT74), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n411), .A2(new_n412), .B1(G33), .B2(G283), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(KEYINPUT74), .A3(new_n416), .A4(new_n418), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n264), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G41), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n251), .A2(G45), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT75), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n429));
  INV_X1    g0229(.A(G45), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(G1), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT5), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G41), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G257), .A3(new_n266), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT77), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT77), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n436), .A2(new_n439), .A3(G257), .A4(new_n266), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT78), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT75), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n432), .B1(new_n431), .B2(new_n434), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT76), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n264), .B1(KEYINPUT5), .B2(new_n425), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n428), .A2(new_n447), .A3(new_n435), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n445), .A2(G274), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n441), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n442), .B1(new_n441), .B2(new_n449), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n275), .B(new_n424), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n341), .A2(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n282), .A2(G77), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT72), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n336), .A2(new_n337), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT6), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT73), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT73), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT6), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n458), .A2(new_n460), .B1(new_n262), .B2(G107), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n262), .A2(G107), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n461), .B(new_n462), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n455), .B1(new_n456), .B2(new_n215), .C1(new_n229), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n453), .B1(new_n464), .B2(new_n281), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n251), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n341), .A2(new_n466), .A3(new_n228), .A4(new_n280), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n262), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n421), .A2(new_n264), .A3(new_n423), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n441), .A2(new_n449), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n441), .A2(new_n442), .A3(new_n449), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n452), .B(new_n468), .C1(new_n473), .C2(G169), .ZN(new_n474));
  OAI211_X1 g0274(.A(G190), .B(new_n424), .C1(new_n450), .C2(new_n451), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n467), .A2(new_n262), .ZN(new_n476));
  AOI211_X1 g0276(.A(new_n453), .B(new_n476), .C1(new_n464), .C2(new_n281), .ZN(new_n477));
  INV_X1    g0277(.A(G200), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n475), .B(new_n477), .C1(new_n473), .C2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n308), .A2(new_n229), .A3(G68), .ZN(new_n480));
  NOR3_X1   g0280(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(G20), .B1(G33), .B2(G97), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT19), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n285), .A2(new_n484), .A3(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT80), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n281), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n368), .A2(new_n370), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n467), .A2(new_n368), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  MUX2_X1   g0295(.A(G238), .B(G244), .S(G1698), .Z(new_n496));
  AOI22_X1  g0296(.A1(new_n308), .A2(new_n496), .B1(G33), .B2(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n266), .ZN(new_n498));
  INV_X1    g0298(.A(G250), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n427), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n431), .A2(new_n253), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n266), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT79), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT79), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n266), .A2(new_n504), .A3(new_n500), .A4(new_n501), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n498), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n275), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n505), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n266), .B2(new_n497), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n272), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n495), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n491), .B(new_n492), .C1(new_n512), .C2(new_n467), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n508), .B(G190), .C1(new_n266), .C2(new_n497), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n506), .B2(new_n478), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n474), .A2(new_n479), .A3(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(G257), .A2(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n216), .A2(G1698), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n308), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n335), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n264), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n436), .A2(G270), .A3(new_n266), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n449), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  OR3_X1    g0327(.A1(new_n467), .A2(KEYINPUT82), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT82), .B1(new_n467), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n417), .B(new_n229), .C1(G33), .C2(new_n262), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(G20), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n281), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n370), .A2(new_n527), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n526), .A2(new_n537), .A3(G169), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT83), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  INV_X1    g0342(.A(new_n537), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n526), .A2(KEYINPUT21), .A3(G169), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n524), .A2(new_n449), .A3(G179), .A4(new_n525), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n306), .A2(new_n307), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT22), .A3(G87), .A4(new_n258), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G116), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n229), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n335), .A2(new_n229), .A3(G87), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n215), .A2(G20), .ZN(new_n556));
  XOR2_X1   g0356(.A(new_n556), .B(KEYINPUT23), .Z(new_n557));
  NAND3_X1  g0357(.A1(new_n552), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n552), .A2(KEYINPUT24), .A3(new_n555), .A4(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n281), .A3(new_n561), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n467), .A2(new_n215), .ZN(new_n563));
  INV_X1    g0363(.A(new_n291), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n556), .ZN(new_n565));
  XOR2_X1   g0365(.A(new_n565), .B(KEYINPUT25), .Z(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G257), .A2(G1698), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n323), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n499), .A2(G1698), .ZN(new_n572));
  XOR2_X1   g0372(.A(KEYINPUT85), .B(G294), .Z(new_n573));
  AOI22_X1  g0373(.A1(new_n308), .A2(new_n572), .B1(new_n573), .B2(G33), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n308), .A2(KEYINPUT84), .A3(G257), .A4(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT86), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n264), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(new_n449), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n436), .A2(G264), .A3(new_n266), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n264), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(KEYINPUT86), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n404), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n576), .B2(new_n264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n449), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n478), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n568), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n272), .B1(new_n579), .B2(new_n582), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n585), .A2(new_n275), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n526), .A2(G200), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n543), .C1(new_n404), .C2(new_n526), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n547), .A2(new_n588), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n410), .A2(new_n518), .A3(new_n595), .ZN(G372));
  INV_X1    g0396(.A(new_n401), .ZN(new_n597));
  INV_X1    g0397(.A(new_n301), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT17), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n353), .B(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n598), .B(new_n600), .C1(new_n298), .C2(new_n373), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n601), .A2(new_n349), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n597), .B1(new_n602), .B2(new_n399), .ZN(new_n603));
  INV_X1    g0403(.A(new_n474), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(KEYINPUT26), .A3(new_n517), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT26), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n474), .B2(new_n516), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n474), .A2(new_n479), .A3(new_n517), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n547), .A2(new_n592), .B1(new_n568), .B2(new_n587), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n611), .A3(new_n511), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n603), .B1(new_n410), .B2(new_n613), .ZN(G369));
  NAND2_X1  g0414(.A1(new_n588), .A2(new_n592), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n544), .A2(new_n545), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n537), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n538), .A2(new_n539), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n620), .A3(new_n540), .ZN(new_n621));
  OR3_X1    g0421(.A1(new_n564), .A2(KEYINPUT27), .A3(G20), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT27), .B1(new_n564), .B2(G20), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(G213), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g0424(.A(KEYINPUT87), .B(G343), .Z(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n615), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n592), .A2(new_n627), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n630), .A2(KEYINPUT88), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT88), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G330), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n617), .A2(new_n620), .A3(new_n540), .A4(new_n594), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n543), .A2(new_n628), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n621), .A2(new_n637), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n568), .A2(new_n628), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n615), .A2(new_n641), .B1(new_n592), .B2(new_n628), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0446(.A(new_n208), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(G41), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n481), .A2(new_n527), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G1), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n233), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT28), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n612), .A2(new_n628), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT29), .ZN(new_n655));
  INV_X1    g0455(.A(new_n511), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n605), .B2(new_n607), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n627), .B1(new_n657), .B2(new_n611), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n424), .B(new_n584), .C1(new_n450), .C2(new_n451), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n545), .A2(new_n509), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n584), .A4(new_n665), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n424), .B1(new_n450), .B2(new_n451), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n526), .A2(new_n275), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n509), .A3(new_n585), .A4(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n627), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n595), .A2(new_n518), .A3(new_n627), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT31), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT90), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n667), .A2(new_n677), .A3(new_n671), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n668), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n667), .B2(new_n671), .ZN(new_n680));
  OAI211_X1 g0480(.A(KEYINPUT31), .B(new_n627), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n635), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n653), .B1(new_n685), .B2(G1), .ZN(G364));
  XOR2_X1   g0486(.A(new_n640), .B(KEYINPUT91), .Z(new_n687));
  NOR2_X1   g0487(.A1(new_n290), .A2(G20), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G45), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n649), .A2(G1), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n638), .A2(new_n639), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n687), .B(new_n690), .C1(G330), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n228), .B1(G20), .B2(new_n272), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(G20), .A2(G179), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n695), .A2(new_n404), .A3(G200), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G322), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n229), .A2(G179), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G190), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G329), .ZN(new_n704));
  INV_X1    g0504(.A(new_n695), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(KEYINPUT95), .A3(G200), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT95), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n695), .B2(new_n478), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G190), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  XOR2_X1   g0511(.A(KEYINPUT33), .B(G317), .Z(new_n712));
  OAI211_X1 g0512(.A(new_n261), .B(new_n704), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n709), .A2(new_n404), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT96), .B(G326), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G283), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n700), .A2(new_n404), .A3(G200), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n404), .A2(G179), .A3(G200), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n229), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n699), .B(new_n719), .C1(new_n573), .C2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n700), .A2(G190), .A3(G200), .ZN(new_n724));
  INV_X1    g0524(.A(G311), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n705), .A2(new_n701), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n723), .B1(new_n522), .B2(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n718), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G107), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n711), .B2(new_n213), .ZN(new_n730));
  INV_X1    g0530(.A(new_n724), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G87), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT32), .ZN(new_n733));
  INV_X1    g0533(.A(G159), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n702), .A2(new_n734), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n732), .B1(new_n204), .B2(new_n726), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n335), .B1(new_n697), .B2(new_n221), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n702), .A2(KEYINPUT32), .A3(new_n734), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n730), .A2(new_n736), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n714), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n739), .B1(new_n219), .B2(new_n740), .C1(new_n262), .C2(new_n721), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n694), .B1(new_n727), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n690), .B(KEYINPUT92), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT94), .Z(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n693), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n246), .A2(G45), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n308), .A2(new_n647), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n751), .B(new_n752), .C1(G45), .C2(new_n233), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n335), .A2(new_n208), .ZN(new_n754));
  INV_X1    g0554(.A(G355), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n755), .B1(G116), .B2(new_n208), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT93), .Z(new_n757));
  AOI21_X1  g0557(.A(new_n750), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n742), .A2(new_n743), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n691), .B2(new_n747), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n692), .A2(new_n760), .ZN(G396));
  INV_X1    g0561(.A(new_n743), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n693), .A2(new_n744), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT97), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n721), .A2(new_n262), .B1(new_n697), .B2(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n765), .A2(new_n767), .B1(new_n714), .B2(G303), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n768), .B1(new_n765), .B2(new_n767), .C1(new_n717), .C2(new_n711), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n718), .A2(new_n512), .B1(new_n702), .B2(new_n725), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n769), .A2(new_n335), .A3(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n771), .B1(new_n215), .B2(new_n724), .C1(new_n527), .C2(new_n726), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n703), .A2(G132), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n718), .A2(new_n213), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n710), .A2(G150), .B1(G143), .B2(new_n696), .ZN(new_n775));
  INV_X1    g0575(.A(G137), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n775), .B1(new_n776), .B2(new_n740), .C1(new_n734), .C2(new_n726), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT34), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n773), .B(new_n774), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n308), .B1(new_n721), .B2(new_n221), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G50), .B2(new_n731), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n781), .C1(new_n778), .C2(new_n777), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT98), .Z(new_n784));
  OAI221_X1 g0584(.A(new_n762), .B1(G77), .B2(new_n764), .C1(new_n784), .C2(new_n694), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n373), .A2(new_n627), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n372), .A2(new_n627), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n408), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(new_n788), .B2(new_n373), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n744), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT99), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n654), .A2(new_n790), .ZN(new_n793));
  INV_X1    g0593(.A(new_n607), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n474), .A2(new_n516), .A3(new_n606), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n511), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n609), .A2(new_n610), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n628), .B(new_n789), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(new_n682), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n690), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n792), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G384));
  INV_X1    g0603(.A(new_n463), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n527), .B1(new_n804), .B2(KEYINPUT35), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n805), .B(new_n230), .C1(KEYINPUT35), .C2(new_n804), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT100), .Z(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT36), .ZN(new_n808));
  OAI21_X1  g0608(.A(G77), .B1(new_n221), .B2(new_n213), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n233), .A2(new_n809), .B1(G50), .B2(new_n213), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(G1), .A3(new_n290), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n297), .B(new_n627), .C1(new_n279), .C2(new_n598), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n297), .A2(new_n627), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n301), .B(new_n813), .C1(new_n376), .C2(new_n296), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n624), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n333), .A2(new_n281), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT16), .B1(new_n327), .B2(new_n332), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n344), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n816), .B(new_n819), .C1(new_n600), .C2(new_n349), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT37), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n346), .A2(new_n347), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n346), .A2(new_n816), .ZN(new_n824));
  AND4_X1   g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n353), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n318), .A2(new_n320), .A3(new_n624), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n822), .B1(new_n827), .B2(new_n353), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n821), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n828), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n823), .A2(new_n824), .A3(new_n822), .A4(new_n353), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(KEYINPUT101), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n820), .A2(new_n829), .A3(new_n832), .A4(KEYINPUT38), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n820), .A2(new_n829), .A3(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n786), .ZN(new_n837));
  AOI221_X4 g0637(.A(new_n815), .B1(new_n833), .B2(new_n836), .C1(new_n798), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n350), .A2(new_n816), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT102), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n815), .B1(new_n798), .B2(new_n837), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n836), .A2(new_n833), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT102), .ZN(new_n844));
  INV_X1    g0644(.A(new_n839), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n836), .A2(KEYINPUT39), .A3(new_n833), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n831), .B(KEYINPUT104), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n823), .A2(KEYINPUT103), .A3(new_n353), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n824), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT103), .B1(new_n823), .B2(new_n353), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n824), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n355), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n833), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n847), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n298), .A2(new_n627), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n840), .A2(new_n846), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n302), .A2(new_n378), .A3(new_n409), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT105), .B1(new_n661), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(KEYINPUT29), .B(new_n627), .C1(new_n657), .C2(new_n611), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n659), .B1(new_n612), .B2(new_n628), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT105), .B(new_n864), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n603), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n863), .B(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n790), .B1(new_n812), .B2(new_n814), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n627), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT106), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n672), .A2(KEYINPUT106), .A3(KEYINPUT31), .A4(new_n627), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n673), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n615), .A2(new_n636), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n609), .A3(new_n628), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(KEYINPUT31), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n842), .B(new_n872), .C1(new_n877), .C2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n875), .A2(new_n876), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n676), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n848), .A2(new_n852), .B1(new_n355), .B2(new_n854), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n833), .B1(new_n887), .B2(KEYINPUT38), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n888), .A4(new_n872), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n886), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n410), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(G330), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n871), .A2(new_n894), .B1(new_n251), .B2(new_n688), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT107), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n871), .A2(new_n894), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT108), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n808), .B(new_n811), .C1(new_n896), .C2(new_n898), .ZN(G367));
  AND2_X1   g0699(.A1(new_n513), .A2(new_n627), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n516), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n656), .A2(new_n900), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT110), .Z(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n604), .A2(new_n627), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n474), .B(new_n479), .C1(new_n477), .C2(new_n628), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n630), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT42), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n474), .B1(new_n909), .B2(new_n592), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n628), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n907), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n643), .A2(new_n911), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n648), .B(KEYINPUT41), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n634), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT44), .B1(new_n925), .B2(new_n910), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT44), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n634), .A2(new_n927), .A3(new_n911), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n910), .B1(new_n632), .B2(new_n633), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT45), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n644), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT45), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n930), .B(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n934), .A2(new_n643), .A3(new_n926), .A4(new_n928), .ZN(new_n935));
  INV_X1    g0735(.A(new_n629), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n630), .B1(new_n642), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n687), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n640), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(new_n937), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n932), .A2(new_n935), .A3(new_n685), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n924), .B1(new_n942), .B2(new_n685), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n689), .A2(G1), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n922), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT111), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n922), .B(KEYINPUT111), .C1(new_n944), .C2(new_n943), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n702), .A2(new_n776), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n711), .A2(new_n734), .B1(new_n388), .B2(new_n697), .ZN(new_n951));
  INV_X1    g0751(.A(new_n726), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n950), .B(new_n951), .C1(G50), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n722), .A2(G68), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n731), .A2(G58), .B1(new_n728), .B2(G77), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n261), .B1(new_n714), .B2(G143), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n718), .A2(new_n262), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n710), .B2(new_n573), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n215), .B2(new_n721), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT112), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n724), .B2(new_n527), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n952), .A2(G283), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n703), .A2(G317), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n963), .A2(new_n961), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n731), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n308), .B1(G303), .B2(new_n696), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n740), .A2(new_n725), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n957), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n693), .ZN(new_n975));
  INV_X1    g0775(.A(new_n752), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n749), .B1(new_n208), .B2(new_n368), .C1(new_n242), .C2(new_n976), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n975), .A2(new_n762), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n905), .A2(new_n747), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n949), .A2(new_n980), .ZN(G387));
  NAND2_X1  g0781(.A1(new_n685), .A2(new_n941), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n649), .B1(new_n684), .B2(new_n940), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n642), .A2(new_n747), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n752), .B1(new_n239), .B2(new_n430), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n650), .B2(new_n754), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n366), .A2(new_n219), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT50), .Z(new_n989));
  NAND2_X1  g0789(.A1(G68), .A2(G77), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n989), .A2(new_n430), .A3(new_n990), .A4(new_n650), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n647), .A2(new_n215), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n750), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n696), .A2(G50), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n388), .B2(new_n702), .C1(new_n711), .C2(new_n343), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n740), .A2(new_n734), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n726), .A2(new_n213), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n996), .A2(new_n958), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n731), .A2(G77), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n721), .A2(new_n368), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n999), .A2(new_n308), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n710), .A2(G311), .B1(G317), .B2(new_n696), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n522), .B2(new_n726), .C1(new_n698), .C2(new_n740), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT48), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n731), .A2(new_n573), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n717), .C2(new_n721), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n728), .A2(G116), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n703), .A2(new_n715), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n323), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1003), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n743), .B(new_n994), .C1(new_n1015), .C2(new_n693), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n941), .A2(new_n944), .B1(new_n985), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n984), .A2(new_n1017), .ZN(G393));
  NAND2_X1  g0818(.A1(new_n932), .A2(new_n935), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n982), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1020), .A2(new_n648), .A3(new_n942), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n932), .A2(new_n944), .A3(new_n935), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n749), .B1(new_n249), .B2(new_n976), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G97), .B2(new_n647), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n714), .A2(G150), .B1(G159), .B2(new_n696), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n711), .A2(new_n219), .B1(new_n512), .B2(new_n718), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n721), .A2(new_n204), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n731), .A2(G68), .B1(new_n952), .B2(new_n366), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n323), .B1(G143), .B2(new_n703), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n714), .A2(G317), .B1(G311), .B2(new_n696), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n261), .B(new_n729), .C1(new_n711), .C2(new_n522), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n724), .A2(new_n717), .B1(new_n702), .B2(new_n698), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT113), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1038), .A2(new_n1039), .B1(new_n722), .B2(G116), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(new_n766), .C2(new_n726), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1033), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n743), .B(new_n1024), .C1(new_n1043), .C2(new_n693), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n910), .B2(new_n747), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1021), .A2(new_n1022), .A3(new_n1045), .ZN(G390));
  AOI21_X1  g0846(.A(new_n786), .B1(new_n658), .B2(new_n789), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n681), .ZN(new_n1048));
  OAI211_X1 g0848(.A(G330), .B(new_n789), .C1(new_n881), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n815), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n635), .B1(new_n676), .B2(new_n885), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n872), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT114), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n815), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1051), .B2(new_n789), .ZN(new_n1056));
  OAI211_X1 g0856(.A(G330), .B(new_n872), .C1(new_n881), .C2(new_n1048), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1047), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1054), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(G330), .B(new_n789), .C1(new_n877), .C2(new_n881), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n815), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1061), .A2(KEYINPUT114), .A3(new_n1047), .A4(new_n1057), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1053), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n892), .A2(G330), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(new_n603), .C1(new_n865), .C2(new_n869), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n888), .B1(new_n298), .B2(new_n627), .C1(new_n1047), .C2(new_n815), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n859), .B1(new_n861), .B2(new_n841), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1057), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1069), .A2(new_n1068), .B1(new_n872), .B2(new_n1051), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1073), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1066), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1076), .A3(new_n648), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n944), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n731), .A2(G150), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT53), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n722), .A2(G159), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n728), .A2(G50), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT54), .B(G143), .Z(new_n1083));
  AOI21_X1  g0883(.A(new_n261), .B1(new_n952), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n714), .A2(G128), .B1(G132), .B2(new_n696), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT115), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(G125), .C2(new_n703), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(KEYINPUT53), .B2(new_n1079), .C1(new_n776), .C2(new_n711), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT116), .Z(new_n1090));
  INV_X1    g0890(.A(KEYINPUT117), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n732), .B2(new_n261), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1029), .B(new_n1092), .C1(G283), .C2(new_n714), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n702), .A2(new_n766), .B1(new_n726), .B2(new_n262), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n774), .B(new_n1094), .C1(G116), .C2(new_n696), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n732), .A2(new_n1091), .A3(new_n261), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G107), .B2(new_n710), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n693), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n743), .B1(new_n343), .B2(new_n763), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n860), .C2(new_n745), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1077), .A2(new_n1078), .A3(new_n1101), .ZN(G378));
  AND3_X1   g0902(.A1(new_n840), .A2(new_n862), .A3(new_n846), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n884), .A2(G330), .A3(new_n889), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n401), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1109), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n399), .A2(new_n401), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n394), .A2(new_n816), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1104), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT120), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n1115), .A3(KEYINPUT120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1125), .A2(new_n884), .A3(G330), .A4(new_n889), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1103), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n863), .A2(new_n1126), .A3(new_n1119), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT121), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT121), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1065), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1073), .B2(new_n1063), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n648), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1132), .B1(new_n1136), .B2(new_n944), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n744), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n954), .B1(new_n368), .B2(new_n726), .C1(new_n740), .C2(new_n527), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n710), .A2(G97), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n728), .A2(G58), .ZN(new_n1142));
  AND4_X1   g0942(.A1(new_n425), .A2(new_n1141), .A3(new_n323), .A4(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1143), .B(new_n1000), .C1(new_n717), .C2(new_n702), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1140), .B(new_n1144), .C1(G107), .C2(new_n696), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT119), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  INV_X1    g0947(.A(G124), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n259), .B1(new_n702), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n714), .A2(G125), .B1(G128), .B2(new_n696), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n731), .A2(new_n1083), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n710), .A2(G132), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n722), .A2(G150), .B1(G137), .B2(new_n952), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(G41), .B(new_n1149), .C1(new_n1154), .C2(KEYINPUT59), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(KEYINPUT59), .B2(new_n1154), .C1(new_n734), .C2(new_n718), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n425), .B1(new_n323), .B2(new_n259), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n219), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT118), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n693), .B1(new_n1147), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n764), .A2(G50), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1139), .A2(new_n690), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1135), .B1(new_n1134), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n1166), .B2(new_n648), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1137), .A2(new_n1167), .ZN(G375));
  NAND2_X1  g0968(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1053), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1065), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1171), .A2(new_n1066), .A3(new_n924), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT122), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1002), .B(new_n261), .C1(new_n204), .C2(new_n718), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n740), .A2(new_n766), .B1(new_n262), .B2(new_n724), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G116), .B2(new_n710), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n215), .B2(new_n726), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1174), .B(new_n1177), .C1(G283), .C2(new_n696), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n522), .B2(new_n702), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n323), .B1(new_n714), .B2(G132), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n1142), .C1(new_n734), .C2(new_n724), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n710), .B2(new_n1083), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n722), .A2(G50), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n703), .A2(G128), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n952), .A2(G150), .B1(G137), .B2(new_n696), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n694), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n743), .B(new_n1187), .C1(new_n213), .C2(new_n763), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n815), .A2(new_n744), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n944), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1063), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1173), .A2(new_n1193), .ZN(G381));
  INV_X1    g0994(.A(G390), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n949), .A2(new_n1195), .A3(new_n980), .ZN(new_n1196));
  OR2_X1    g0996(.A1(G393), .A2(G396), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1196), .A2(G381), .A3(G384), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(G407));
  NAND2_X1  g1003(.A1(new_n626), .A2(G213), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT124), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1206), .A2(KEYINPUT124), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(G407), .A2(G213), .A3(new_n1207), .A4(new_n1208), .ZN(G409));
  XOR2_X1   g1009(.A(G393), .B(G396), .Z(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G387), .A2(G390), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1196), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1195), .B1(new_n949), .B2(new_n980), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n980), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1215), .B(G390), .C1(new_n947), .C2(new_n948), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1214), .A2(new_n1216), .A3(new_n1210), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1164), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1127), .B(new_n863), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n1191), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1134), .A2(new_n923), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1221), .B1(new_n1132), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT125), .B1(new_n1224), .B2(G378), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1137), .A2(G378), .A3(new_n1167), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1078), .A2(new_n1101), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n649), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n1076), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1222), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1229), .B(new_n1230), .C1(new_n1231), .C2(new_n1221), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1225), .A2(new_n1226), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT60), .B1(new_n1171), .B2(new_n1066), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n649), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G384), .B1(new_n1238), .B2(new_n1193), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n802), .B(new_n1192), .C1(new_n1234), .C2(new_n1237), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1233), .A2(KEYINPUT63), .A3(new_n1204), .A4(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1218), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1233), .A2(new_n1204), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1239), .A2(new_n1240), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1205), .A2(G2897), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1246), .B(new_n1249), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1247), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1245), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1254), .A2(KEYINPUT63), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1233), .A2(new_n1204), .A3(new_n1241), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1243), .B(new_n1244), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT127), .B1(new_n1254), .B2(new_n1244), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT127), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1260), .B(KEYINPUT61), .C1(new_n1245), .C2(new_n1253), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1233), .A2(new_n1263), .A3(new_n1204), .A4(new_n1241), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1259), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1258), .B1(new_n1266), .B2(new_n1218), .ZN(G405));
  NAND2_X1  g1067(.A1(G375), .A2(new_n1229), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1226), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1218), .B(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1241), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1218), .A2(new_n1269), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1218), .A2(new_n1269), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1241), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(G402));
endmodule


