//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT71), .ZN(new_n204));
  INV_X1    g003(.A(G15gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G43gat), .ZN(new_n207));
  XOR2_X1   g006(.A(G183gat), .B(G190gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT24), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT24), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT23), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n218), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n212), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n212), .A2(new_n223), .A3(new_n225), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT64), .B(G176gat), .Z(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT23), .A3(new_n214), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n214), .A2(new_n215), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(new_n216), .B2(new_n217), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n229), .A2(new_n209), .A3(new_n211), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n213), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n237), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n219), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n210), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n236), .B2(new_n235), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n238), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(KEYINPUT1), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT69), .B(G113gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(G120gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT68), .B(G120gat), .Z(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n251), .B1(new_n250), .B2(G120gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G113gat), .B2(G120gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n248), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n224), .A2(new_n225), .B1(new_n213), .B2(new_n232), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n245), .B1(new_n264), .B2(new_n227), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(G227gat), .A2(G233gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT33), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n207), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(KEYINPUT32), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n268), .B1(new_n263), .B2(new_n267), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275));
  OR3_X1    g074(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT34), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT34), .B1(new_n274), .B2(new_n275), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n269), .B(KEYINPUT32), .C1(new_n270), .C2(new_n207), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n273), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n273), .A2(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n202), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n277), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT36), .A3(new_n279), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G148gat), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n288), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT81), .B1(new_n288), .B2(G141gat), .ZN(new_n290));
  INV_X1    g089(.A(G141gat), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(G148gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n292), .A2(new_n293), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n295), .A2(KEYINPUT78), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(KEYINPUT78), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n302), .A2(new_n303), .B1(new_n297), .B2(new_n298), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n295), .B1(new_n305), .B2(KEYINPUT2), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n296), .A2(KEYINPUT79), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n288), .A2(G141gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n291), .A2(G148gat), .ZN(new_n309));
  OAI22_X1  g108(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(KEYINPUT80), .A3(new_n310), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n301), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n266), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n315), .A2(new_n313), .B1(new_n294), .B2(new_n300), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n262), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT85), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT84), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT85), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n324), .A3(new_n266), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT5), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n301), .B(new_n328), .C1(new_n314), .C2(new_n316), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n329), .B(new_n266), .C1(new_n319), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n320), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n323), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n262), .A2(new_n319), .A3(KEYINPUT4), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n331), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT0), .ZN(new_n342));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n346));
  INV_X1    g145(.A(new_n344), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n337), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n348), .A2(new_n346), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI211_X1 g156(.A(new_n245), .B(new_n357), .C1(new_n264), .C2(new_n227), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n234), .B2(new_n246), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT22), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(KEYINPUT73), .B1(G211gat), .B2(G218gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(KEYINPUT73), .B2(new_n361), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n365), .A2(KEYINPUT74), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(new_n364), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI22_X1  g170(.A1(new_n358), .A2(new_n360), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n234), .A2(new_n246), .A3(new_n356), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n368), .A2(new_n371), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n373), .B(new_n374), .C1(new_n265), .C2(new_n359), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n372), .A2(KEYINPUT75), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n358), .A2(new_n360), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n374), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n355), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n376), .B2(new_n379), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n385), .A2(new_n386), .A3(new_n354), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n380), .A2(KEYINPUT30), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT77), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n386), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n355), .A3(new_n384), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n388), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n382), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G22gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n374), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n319), .B1(new_n400), .B2(new_n330), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n374), .B1(new_n329), .B2(new_n399), .ZN(new_n402));
  OAI211_X1 g201(.A(G228gat), .B(G233gat), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n369), .A2(KEYINPUT86), .A3(new_n366), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n366), .B(KEYINPUT86), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n399), .C1(new_n369), .C2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n407), .A2(new_n328), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n408), .B2(new_n319), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n409), .A2(new_n402), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT31), .B(G50gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n403), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n403), .B2(new_n410), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n398), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n403), .A2(new_n410), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n411), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(new_n397), .A3(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n287), .B1(new_n395), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n348), .A2(KEYINPUT87), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n321), .A2(new_n325), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n334), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n323), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n427), .A3(KEYINPUT39), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n344), .B1(new_n427), .B2(KEYINPUT39), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n427), .A2(KEYINPUT39), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n432), .A2(KEYINPUT40), .A3(new_n428), .A4(new_n344), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n337), .A2(new_n339), .A3(new_n434), .A4(new_n347), .ZN(new_n435));
  AND4_X1   g234(.A1(new_n422), .A2(new_n431), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n381), .A2(new_n351), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n392), .A2(new_n388), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n420), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT6), .B1(new_n340), .B2(new_n344), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(new_n422), .A3(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n440), .A2(new_n422), .A3(KEYINPUT88), .A4(new_n435), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n350), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n385), .A2(new_n386), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n376), .A2(new_n379), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n354), .B1(new_n448), .B2(new_n446), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT38), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n372), .A2(new_n375), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT38), .B1(new_n452), .B2(KEYINPUT37), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n380), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n439), .B1(new_n445), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n420), .B1(new_n285), .B2(new_n279), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n382), .A2(new_n390), .A3(new_n457), .A4(new_n394), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n416), .A2(new_n419), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n460), .B(new_n461), .C1(new_n280), .C2(new_n281), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n438), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n445), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n421), .A2(new_n456), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT15), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  INV_X1    g266(.A(G50gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(G43gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(G43gat), .ZN(new_n470));
  INV_X1    g269(.A(G43gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(G50gat), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n466), .B(new_n469), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G29gat), .ZN(new_n474));
  INV_X1    g273(.A(G36gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n474), .A3(new_n475), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT14), .A3(new_n477), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n471), .A2(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n468), .A2(G43gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n484), .B(new_n485), .C1(new_n467), .C2(KEYINPUT15), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n473), .A2(new_n480), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n470), .A2(new_n472), .A3(new_n466), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n477), .A2(KEYINPUT14), .ZN(new_n489));
  NOR3_X1   g288(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n477), .A2(KEYINPUT14), .B1(new_n474), .B2(new_n475), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT91), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n487), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499));
  INV_X1    g298(.A(G1gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT16), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(G1gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n502), .A2(new_n503), .A3(G8gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n498), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n510), .A3(new_n497), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n495), .A2(new_n513), .A3(new_n510), .A4(new_n497), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n508), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n494), .A2(new_n510), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n509), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  AOI211_X1 g319(.A(KEYINPUT94), .B(KEYINPUT18), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n487), .A2(new_n496), .A3(new_n493), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n496), .B1(new_n487), .B2(new_n493), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n513), .B1(new_n525), .B2(new_n510), .ZN(new_n526));
  INV_X1    g325(.A(new_n514), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n509), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n520), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n522), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n521), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(KEYINPUT18), .A3(new_n520), .A4(new_n529), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n498), .B2(new_n508), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n520), .B(KEYINPUT13), .Z(new_n538));
  NAND3_X1  g337(.A1(new_n516), .A2(new_n525), .A3(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G197gat), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT11), .B(G169gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT12), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n534), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n531), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(new_n540), .A3(new_n534), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n533), .A2(new_n547), .B1(new_n549), .B2(new_n545), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n297), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G64gat), .Z(new_n555));
  INV_X1    g354(.A(G71gat), .ZN(new_n556));
  INV_X1    g355(.A(G78gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n559), .B(new_n558), .C1(new_n564), .C2(new_n561), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT95), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT95), .B1(new_n563), .B2(new_n565), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n554), .B1(new_n569), .B2(new_n508), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n554), .A3(new_n508), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n553), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n574), .A2(new_n570), .A3(new_n552), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n563), .A2(new_n565), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n568), .ZN(new_n578));
  AND2_X1   g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G127gat), .ZN(new_n583));
  INV_X1    g382(.A(G127gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n583), .B2(new_n585), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n576), .A2(new_n590), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n573), .A2(new_n575), .B1(new_n588), .B2(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G120gat), .B(G148gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT103), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(G85gat), .B(G92gat), .C1(KEYINPUT97), .C2(KEYINPUT7), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n605), .B(new_n607), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT8), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT98), .B1(G99gat), .B2(G106gat), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n602), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n615), .B1(new_n612), .B2(new_n613), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n613), .B2(new_n612), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n610), .A2(new_n609), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n606), .B1(new_n604), .B2(new_n603), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n601), .A4(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(KEYINPUT99), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n611), .A2(new_n617), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n601), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n577), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n618), .A2(new_n623), .A3(new_n565), .A4(new_n563), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n566), .A2(new_n567), .A3(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n600), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n599), .B1(new_n628), .B2(new_n629), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n598), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(KEYINPUT104), .B(new_n598), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT102), .B1(new_n631), .B2(new_n634), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n631), .A2(KEYINPUT102), .A3(new_n634), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n599), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n636), .A2(new_n598), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n495), .A3(new_n497), .ZN(new_n651));
  NAND3_X1  g450(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n651), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT100), .B1(new_n651), .B2(new_n652), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n633), .A2(new_n517), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n512), .B2(new_n514), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n650), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G134gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n298), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n515), .A2(new_n656), .ZN(new_n665));
  INV_X1    g464(.A(new_n650), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n665), .B(new_n666), .C1(new_n653), .C2(new_n654), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n661), .A2(new_n664), .B1(new_n659), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n659), .A2(new_n667), .A3(KEYINPUT101), .A4(new_n664), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n594), .B(new_n649), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n465), .A2(new_n550), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n349), .A2(new_n350), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n672), .A2(new_n438), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n672), .A2(new_n438), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G8gat), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n681), .B2(new_n679), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n689), .B(KEYINPUT106), .C1(new_n683), .C2(new_n682), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1325gat));
  NOR2_X1   g490(.A1(new_n280), .A2(new_n281), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n672), .A2(new_n205), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n672), .A2(new_n287), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n205), .ZN(G1326gat));
  NAND2_X1  g495(.A1(new_n672), .A2(new_n420), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT107), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n421), .A2(new_n456), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n459), .A2(new_n464), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n548), .A2(KEYINPUT94), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n530), .A2(new_n522), .A3(new_n531), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n547), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n549), .A2(new_n545), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n594), .A2(new_n648), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n659), .A2(new_n667), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n665), .B1(new_n653), .B2(new_n654), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT101), .B1(new_n712), .B2(new_n650), .ZN(new_n713));
  INV_X1    g512(.A(new_n664), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n669), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n703), .A2(new_n708), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n474), .A3(new_n674), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n465), .B2(new_n716), .ZN(new_n723));
  INV_X1    g522(.A(new_n716), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n550), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n673), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n721), .A2(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(new_n438), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n718), .A2(new_n475), .A3(new_n438), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(KEYINPUT109), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(KEYINPUT109), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n732), .B(new_n737), .C1(new_n735), .C2(new_n733), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n725), .A3(new_n287), .A4(new_n727), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n692), .A2(G43gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n703), .A2(new_n741), .A3(new_n708), .A4(new_n717), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n742), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT47), .B1(new_n745), .B2(new_n740), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI211_X1 g547(.A(KEYINPUT111), .B(KEYINPUT47), .C1(new_n745), .C2(new_n740), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(G1330gat));
  NAND4_X1  g549(.A1(new_n723), .A2(new_n725), .A3(new_n420), .A4(new_n727), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n718), .A2(new_n468), .A3(new_n420), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT48), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n754), .B(new_n756), .ZN(G1331gat));
  AOI21_X1  g556(.A(new_n593), .B1(new_n715), .B2(new_n669), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n758), .A2(new_n550), .A3(new_n648), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n703), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n703), .A2(KEYINPUT113), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n674), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g566(.A1(new_n764), .A2(new_n731), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  INV_X1    g571(.A(new_n287), .ZN(new_n773));
  OAI21_X1  g572(.A(G71gat), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n693), .A2(new_n556), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n764), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1334gat));
  NOR2_X1   g577(.A1(new_n764), .A2(new_n460), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n557), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n465), .A2(new_n716), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n708), .A2(new_n594), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT51), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  INV_X1    g583(.A(new_n782), .ZN(new_n785));
  NOR4_X1   g584(.A1(new_n465), .A2(new_n784), .A3(new_n716), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OR4_X1    g586(.A1(G85gat), .A2(new_n787), .A3(new_n673), .A4(new_n649), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n785), .A2(new_n649), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n726), .A2(new_n674), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G85gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n465), .A2(new_n716), .A3(new_n785), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n784), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(G92gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n438), .A2(new_n799), .A3(new_n648), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT115), .Z(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n703), .A2(new_n724), .A3(new_n782), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n726), .A2(new_n789), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n731), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n807), .B2(new_n799), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI221_X1 g609(.A(new_n810), .B1(new_n787), .B2(new_n801), .C1(new_n807), .C2(new_n799), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1337gat));
  OR4_X1    g611(.A1(G99gat), .A2(new_n787), .A3(new_n692), .A4(new_n649), .ZN(new_n813));
  OAI21_X1  g612(.A(G99gat), .B1(new_n806), .B2(new_n773), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1338gat));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n460), .A2(G106gat), .A3(new_n649), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n783), .B2(new_n786), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n723), .A2(new_n725), .A3(new_n420), .A4(new_n789), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n798), .A2(new_n804), .A3(new_n817), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n820), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n816), .B(new_n822), .C1(new_n824), .C2(new_n821), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n821), .B1(new_n823), .B2(new_n820), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1339gat));
  AND2_X1   g628(.A1(new_n537), .A2(new_n539), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n830), .A2(new_n538), .B1(new_n519), .B2(new_n520), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n544), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n706), .A2(new_n648), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n599), .B1(new_n632), .B2(new_n633), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n631), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n835), .B2(new_n631), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n834), .B1(new_n840), .B2(new_n645), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT54), .B(new_n600), .C1(new_n631), .C2(new_n634), .ZN(new_n842));
  INV_X1    g641(.A(new_n598), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT120), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n631), .A2(new_n634), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n599), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n848), .A3(new_n598), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n841), .A2(new_n850), .B1(new_n645), .B2(new_n646), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n842), .A2(KEYINPUT120), .A3(new_n843), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n848), .B1(new_n847), .B2(new_n598), .ZN(new_n853));
  INV_X1    g652(.A(new_n644), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n642), .A3(new_n600), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n631), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT119), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n834), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n833), .B1(new_n550), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n716), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n706), .A2(new_n832), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n864), .A2(new_n861), .A3(new_n716), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n594), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT118), .B1(new_n671), .B2(new_n708), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n758), .A2(new_n550), .A3(new_n868), .A4(new_n649), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT121), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n708), .A2(new_n860), .A3(new_n851), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n724), .B1(new_n872), .B2(new_n833), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n864), .A2(new_n861), .A3(new_n716), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n593), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n867), .A2(new_n869), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n673), .ZN(new_n880));
  INV_X1    g679(.A(new_n457), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n438), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n250), .A3(new_n708), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n731), .A2(new_n674), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n879), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n888), .A2(new_n708), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n890), .B2(new_n253), .ZN(G1340gat));
  NAND3_X1  g690(.A1(new_n888), .A2(new_n648), .A3(new_n889), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G120gat), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n649), .A2(new_n254), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n883), .B2(new_n894), .ZN(G1341gat));
  NAND3_X1  g694(.A1(new_n884), .A2(new_n584), .A3(new_n594), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n888), .A2(new_n594), .A3(new_n889), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n584), .ZN(G1342gat));
  INV_X1    g697(.A(G134gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n724), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT56), .B1(new_n883), .B2(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n883), .A2(KEYINPUT56), .A3(new_n900), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n888), .A2(new_n724), .A3(new_n889), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n899), .ZN(G1343gat));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n287), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n871), .A2(new_n878), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n906), .B2(new_n420), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n420), .A2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n875), .B2(new_n877), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n708), .B(new_n905), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G141gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n287), .A2(new_n460), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n674), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n438), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n550), .A2(G141gat), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n906), .A2(KEYINPUT123), .A3(new_n674), .A4(new_n914), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n912), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  NOR4_X1   g720(.A1(new_n915), .A2(G141gat), .A3(new_n438), .A4(new_n550), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n913), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n912), .A2(new_n913), .A3(new_n920), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n922), .B1(new_n911), .B2(G141gat), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n926), .B(new_n927), .C1(new_n913), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(G1344gat));
  OAI21_X1  g729(.A(new_n875), .B1(new_n708), .B2(new_n671), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n420), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n879), .A2(new_n909), .B1(new_n932), .B2(KEYINPUT57), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n886), .A2(new_n287), .A3(new_n649), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n288), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n907), .A2(new_n910), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n934), .A2(new_n936), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n935), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n917), .A2(new_n919), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n936), .B1(new_n941), .B2(new_n648), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g742(.A(G155gat), .B1(new_n941), .B2(new_n594), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n938), .A2(new_n905), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n593), .A2(new_n297), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT125), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(G1346gat));
  AOI21_X1  g747(.A(G162gat), .B1(new_n941), .B2(new_n724), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n716), .A2(new_n298), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n945), .B2(new_n950), .ZN(G1347gat));
  NAND2_X1  g750(.A1(new_n438), .A2(new_n673), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n879), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n457), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n550), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(new_n214), .ZN(G1348gat));
  NAND4_X1  g755(.A1(new_n953), .A2(new_n693), .A3(new_n460), .A4(new_n648), .ZN(new_n957));
  MUX2_X1   g756(.A(new_n228), .B(G176gat), .S(new_n957), .Z(G1349gat));
  OR3_X1    g757(.A1(new_n954), .A2(new_n235), .A3(new_n593), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n960));
  INV_X1    g759(.A(G183gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n961), .B1(new_n954), .B2(new_n593), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n960), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1350gat));
  OAI22_X1  g764(.A1(new_n954), .A2(new_n716), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(G1351gat));
  NAND4_X1  g767(.A1(new_n933), .A2(new_n673), .A3(new_n438), .A4(new_n773), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(new_n550), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n914), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n708), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n971), .A2(new_n974), .ZN(G1352gat));
  NOR3_X1   g774(.A1(new_n972), .A2(G204gat), .A3(new_n649), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(G204gat), .B1(new_n969), .B2(new_n649), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n977), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(G1353gat));
  NOR3_X1   g780(.A1(new_n972), .A2(G211gat), .A3(new_n593), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n982), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n986), .B1(new_n969), .B2(new_n593), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n988));
  NAND2_X1  g787(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n989), .B(new_n986), .C1(new_n969), .C2(new_n593), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n984), .A2(new_n988), .A3(new_n990), .ZN(G1354gat));
  OAI21_X1  g790(.A(G218gat), .B1(new_n969), .B2(new_n716), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n716), .A2(G218gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(new_n972), .B2(new_n993), .ZN(G1355gat));
endmodule


