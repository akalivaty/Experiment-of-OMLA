//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n482), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n477), .B1(new_n483), .B2(new_n462), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n476), .A2(new_n484), .ZN(G160));
  NOR2_X1   g060(.A1(new_n478), .A2(new_n462), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n478), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G138), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(new_n495), .B1(new_n488), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n472), .A2(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n462), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n463), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G102), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n472), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n506));
  OAI211_X1 g081(.A(KEYINPUT70), .B(new_n503), .C1(new_n506), .C2(new_n462), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n497), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT71), .B(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI211_X1 g090(.A(G50), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G75), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g097(.A(G88), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(G62), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n518), .A2(new_n525), .ZN(G166));
  OAI211_X1 g101(.A(G543), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT72), .B(G51), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT6), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(new_n513), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT5), .B(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT73), .B(KEYINPUT74), .Z(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND4_X1  g120(.A1(new_n534), .A2(G90), .A3(new_n513), .A4(new_n538), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n534), .A2(G52), .A3(G543), .A4(new_n513), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n519), .A2(new_n521), .A3(G64), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(new_n514), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n546), .A2(new_n547), .A3(new_n551), .A4(KEYINPUT75), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(G171));
  NAND4_X1  g131(.A1(new_n534), .A2(G43), .A3(G543), .A4(new_n513), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT76), .B(G81), .Z(new_n558));
  NAND4_X1  g133(.A1(new_n534), .A2(new_n513), .A3(new_n538), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n519), .A2(new_n521), .A3(G56), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n514), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G188));
  NAND3_X1  g147(.A1(new_n519), .A2(new_n521), .A3(G65), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT78), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n573), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(G651), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n513), .B(new_n538), .C1(new_n514), .C2(new_n515), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G91), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(G53), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n527), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n531), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n512), .B1(new_n588), .B2(KEYINPUT6), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n589), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n579), .A2(new_n582), .A3(new_n585), .A4(new_n590), .ZN(G299));
  AND2_X1   g166(.A1(new_n554), .A2(new_n555), .ZN(G301));
  OR2_X1    g167(.A1(new_n518), .A2(new_n525), .ZN(G303));
  NAND3_X1  g168(.A1(new_n589), .A2(G49), .A3(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n534), .A2(G87), .A3(new_n513), .A4(new_n538), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND3_X1  g172(.A1(new_n589), .A2(G86), .A3(new_n538), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n515), .B1(new_n586), .B2(new_n587), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n599), .A2(new_n510), .A3(new_n512), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G48), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n538), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NOR3_X1   g178(.A1(new_n602), .A2(new_n603), .A3(new_n588), .ZN(new_n604));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n522), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT79), .B1(new_n607), .B2(new_n514), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n598), .B(new_n601), .C1(new_n604), .C2(new_n608), .ZN(G305));
  NAND3_X1  g184(.A1(new_n589), .A2(G85), .A3(new_n538), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n589), .A2(G47), .A3(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n522), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n514), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(G290));
  AOI22_X1  g191(.A1(new_n538), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(new_n511), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n600), .A2(G54), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n580), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n589), .A2(G92), .A3(new_n538), .A4(new_n620), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n618), .A2(new_n619), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G171), .B2(new_n626), .ZN(G284));
  OAI21_X1  g203(.A(new_n627), .B1(G171), .B2(new_n626), .ZN(G321));
  NAND2_X1  g204(.A1(G299), .A2(new_n626), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G168), .B2(new_n626), .ZN(G280));
  XNOR2_X1  g206(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g207(.A(new_n625), .ZN(new_n633));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n564), .A2(new_n626), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n625), .A2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n482), .A2(new_n502), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n486), .A2(G123), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n488), .A2(G135), .ZN(new_n647));
  NOR2_X1   g222(.A1(G99), .A2(G2105), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT84), .B(G2096), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2435), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2438), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT14), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n672), .B2(new_n673), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n675), .B1(new_n674), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n681), .B(new_n684), .Z(G227));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n696), .B(new_n697), .C1(new_n695), .C2(new_n694), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(G1986), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G1981), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G35), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT29), .Z(new_n709));
  INV_X1    g284(.A(G2090), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT95), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT31), .B(G11), .Z(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n706), .A2(G26), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n486), .A2(G128), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n488), .A2(G140), .ZN(new_n717));
  NOR2_X1   g292(.A1(G104), .A2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n715), .B1(new_n720), .B2(G29), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n715), .B(new_n721), .S(KEYINPUT28), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2067), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT30), .B(G28), .Z(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(G29), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n488), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n486), .A2(G129), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n502), .A2(G105), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  NAND4_X1  g305(.A1(new_n726), .A2(new_n727), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G32), .B(new_n731), .S(G29), .Z(new_n732));
  XOR2_X1   g307(.A(KEYINPUT27), .B(G1996), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n650), .A2(new_n706), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n706), .A2(G27), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G164), .B2(new_n706), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G2078), .ZN(new_n738));
  NOR4_X1   g313(.A1(new_n725), .A2(new_n734), .A3(new_n735), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G168), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n709), .A2(new_n710), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n565), .B2(new_n746), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1341), .Z(new_n749));
  OR2_X1    g324(.A1(new_n737), .A2(G2078), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n744), .A2(new_n745), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(G299), .A2(G16), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n746), .A2(KEYINPUT23), .A3(G20), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n754));
  INV_X1    g329(.A(G20), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G16), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1956), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n706), .A2(G33), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n488), .A2(G139), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n502), .A2(G103), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n482), .A2(G127), .ZN(new_n763));
  INV_X1    g338(.A(G115), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n463), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n760), .B(new_n762), .C1(new_n765), .C2(G2105), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n706), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2072), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n751), .A2(new_n758), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n714), .A2(new_n739), .A3(new_n743), .A4(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT36), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G24), .ZN(new_n773));
  XOR2_X1   g348(.A(G290), .B(KEYINPUT89), .Z(new_n774));
  AOI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1986), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n706), .A2(G25), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n486), .A2(G119), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n488), .A2(G131), .ZN(new_n780));
  OR2_X1    g355(.A1(G95), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(new_n706), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT35), .B(G1991), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n785), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n746), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n746), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT90), .B(G1971), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G6), .B(G305), .S(G16), .Z(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G16), .B2(G23), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  INV_X1    g374(.A(G1976), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n798), .A2(KEYINPUT33), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(KEYINPUT33), .ZN(new_n803));
  AOI21_X1  g378(.A(G1976), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n792), .B(new_n795), .C1(new_n801), .C2(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n777), .B(new_n788), .C1(new_n805), .C2(KEYINPUT34), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n772), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n771), .A2(KEYINPUT36), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT92), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n772), .B(new_n810), .C1(new_n806), .C2(new_n807), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n770), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G160), .A2(new_n706), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT24), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(G34), .ZN(new_n818));
  AOI21_X1  g393(.A(G29), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n815), .A2(new_n819), .B1(KEYINPUT94), .B2(G2084), .ZN(new_n820));
  NAND2_X1  g395(.A1(KEYINPUT94), .A2(G2084), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  NOR2_X1   g397(.A1(G5), .A2(G16), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G171), .B2(G16), .ZN(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G4), .A2(G16), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n633), .B2(G16), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT93), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n814), .A2(new_n822), .A3(new_n826), .A4(new_n831), .ZN(G150));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g408(.A1(G150), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n831), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n835), .B(new_n770), .C1(new_n812), .C2(new_n813), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n836), .A2(KEYINPUT96), .A3(new_n822), .A4(new_n826), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(G311));
  NAND4_X1  g413(.A1(new_n534), .A2(G93), .A3(new_n513), .A4(new_n538), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n534), .A2(G55), .A3(G543), .A4(new_n513), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n519), .A2(new_n521), .A3(G67), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n514), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT97), .B(G860), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  AOI21_X1  g423(.A(new_n588), .B1(new_n560), .B2(new_n561), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n600), .B2(G43), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n850), .A3(new_n559), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n588), .B1(new_n841), .B2(new_n842), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n600), .B2(G55), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n564), .A2(new_n853), .A3(new_n839), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n633), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n848), .B1(new_n859), .B2(new_n846), .ZN(G145));
  XNOR2_X1  g435(.A(new_n720), .B(new_n731), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n501), .A2(new_n504), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n497), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n766), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  AOI22_X1  g442(.A1(G130), .A2(new_n486), .B1(new_n488), .B2(G142), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT98), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n870), .B(new_n871), .C1(G118), .C2(new_n462), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n783), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n642), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(new_n867), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n650), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G160), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n865), .B(new_n875), .Z(new_n879));
  OAI211_X1 g454(.A(new_n876), .B(new_n878), .C1(new_n879), .C2(new_n867), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n880), .B(new_n881), .C1(new_n879), .C2(new_n878), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n845), .A2(G868), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n796), .A2(G290), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n600), .A2(G47), .B1(new_n514), .B2(new_n614), .ZN(new_n889));
  NAND3_X1  g464(.A1(G288), .A2(new_n889), .A3(new_n610), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(G303), .A2(G305), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n603), .B1(new_n602), .B2(new_n588), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n607), .A2(KEYINPUT79), .A3(new_n514), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n894), .A2(new_n895), .B1(G48), .B2(new_n600), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(G166), .A3(new_n598), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n888), .B1(new_n887), .B2(new_n890), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n892), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n887), .A2(new_n890), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n898), .A2(KEYINPUT102), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT42), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT103), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n855), .B(KEYINPUT100), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n637), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n908));
  NAND2_X1  g483(.A1(G299), .A2(new_n625), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(G299), .A2(new_n625), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(G299), .A2(new_n625), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(KEYINPUT101), .A3(new_n909), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n907), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n910), .B2(new_n911), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n907), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n905), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n904), .A2(KEYINPUT103), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n884), .B(new_n886), .C1(new_n924), .C2(new_n626), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n626), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT104), .B1(new_n926), .B2(new_n885), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(G295));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n885), .ZN(G331));
  NAND3_X1  g504(.A1(G171), .A2(new_n851), .A3(new_n854), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G171), .B1(new_n851), .B2(new_n854), .ZN(new_n932));
  OAI21_X1  g507(.A(G286), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G301), .A2(new_n855), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(G168), .A3(new_n930), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n933), .A2(new_n917), .A3(new_n918), .A4(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n910), .A2(new_n911), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n934), .A2(G168), .A3(new_n930), .ZN(new_n938));
  AOI21_X1  g513(.A(G168), .B1(new_n934), .B2(new_n930), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n940), .A3(new_n903), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n881), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n912), .A2(new_n914), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n938), .B2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n900), .B2(new_n902), .ZN(new_n946));
  INV_X1    g521(.A(new_n899), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n947), .A2(new_n891), .A3(new_n893), .A4(new_n897), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n898), .A2(KEYINPUT102), .A3(new_n901), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT105), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n936), .A2(new_n944), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n942), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n936), .A2(new_n944), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n881), .A4(new_n941), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n936), .A2(new_n940), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n954), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n881), .A4(new_n941), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n958), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n955), .A2(new_n961), .A3(new_n881), .A4(new_n941), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n942), .B1(new_n959), .B2(new_n954), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n961), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n967), .A2(new_n972), .A3(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n863), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n476), .A2(new_n484), .A3(G40), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n720), .B(G2067), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT110), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n731), .B(G1996), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n784), .A2(new_n787), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n783), .A2(new_n786), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G290), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n776), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT109), .Z(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n776), .B2(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n983), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n476), .A2(new_n484), .A3(G40), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n981), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n742), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n508), .A2(new_n978), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g579(.A(G2084), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n497), .B2(new_n862), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n999), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n998), .B1(new_n1010), .B2(G286), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(G168), .A3(new_n1009), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n998), .B1(new_n1012), .B2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n981), .A2(G40), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n471), .A2(new_n475), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n980), .B(G1384), .C1(new_n497), .C2(new_n862), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2078), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1004), .A2(new_n999), .A3(new_n1008), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(new_n825), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT123), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(KEYINPUT123), .ZN(new_n1028));
  XNOR2_X1  g603(.A(G301), .B(KEYINPUT54), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n508), .B2(new_n978), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1030), .A2(new_n982), .A3(new_n1019), .ZN(new_n1031));
  INV_X1    g606(.A(G2078), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT53), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR4_X1   g608(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1016), .B1(new_n1023), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1006), .A2(G40), .A3(new_n476), .A4(new_n484), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n796), .A2(G1976), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT112), .B(G86), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n581), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n896), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n601), .B1(new_n604), .B2(new_n608), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1044), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n896), .A2(new_n1042), .A3(new_n598), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1046), .A2(new_n1051), .A3(G8), .A4(new_n1036), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n800), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1036), .A2(G8), .A3(new_n1037), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1039), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT115), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1039), .A2(new_n1052), .A3(new_n1057), .A4(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1031), .B2(G1971), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1004), .A2(new_n710), .A3(new_n999), .A4(new_n1008), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1003), .A2(new_n980), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(new_n1020), .A3(new_n999), .ZN(new_n1064));
  INV_X1    g639(.A(G1971), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(KEYINPUT111), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n1068), .B(KEYINPUT55), .Z(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(G8), .A3(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1059), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1001), .A2(new_n1021), .A3(G2078), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1025), .A2(new_n1072), .A3(new_n1033), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1029), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1069), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n508), .A2(new_n1007), .A3(new_n978), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n999), .A3(new_n710), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(new_n1080), .C1(new_n1031), .C2(G1971), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1080), .B1(new_n1083), .B2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1076), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1035), .A2(new_n1071), .A3(new_n1075), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n999), .A2(KEYINPUT118), .A3(new_n1006), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1036), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT121), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1095), .B(new_n1092), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1064), .A2(G1996), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1087), .B1(new_n1098), .B2(new_n564), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1077), .A2(new_n999), .A3(new_n1078), .ZN(new_n1101));
  INV_X1    g676(.A(G1956), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1031), .A2(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(KEYINPUT119), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1103), .A2(new_n1107), .A3(KEYINPUT120), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1063), .A2(new_n1020), .A3(new_n999), .A4(new_n1100), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G299), .B(KEYINPUT57), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT119), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(KEYINPUT61), .B(new_n1106), .C1(new_n1108), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT61), .B1(new_n1106), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1095), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1097), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1091), .A2(KEYINPUT121), .A3(new_n1093), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .A3(new_n565), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1099), .A2(new_n1116), .A3(new_n1119), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1091), .A2(G2067), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1024), .A2(new_n830), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(KEYINPUT60), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(new_n633), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(KEYINPUT60), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT120), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1112), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1118), .B1(new_n1138), .B2(KEYINPUT61), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(KEYINPUT122), .A3(new_n1099), .A4(new_n1125), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1133), .A2(new_n625), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1106), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1086), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1067), .A2(G8), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1076), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1010), .A2(G8), .A3(G168), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT116), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1055), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(new_n1148), .A3(new_n1076), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1151), .B(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1085), .A2(new_n1059), .A3(new_n1070), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1145), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1052), .A2(new_n800), .A3(new_n796), .ZN(new_n1160));
  OAI211_X1 g735(.A(G8), .B(new_n1036), .C1(new_n1160), .C2(new_n1041), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1070), .B2(new_n1055), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT113), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1161), .B(KEYINPUT113), .C1(new_n1070), .C2(new_n1055), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1155), .A2(new_n1159), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1158), .A2(G301), .A3(new_n1073), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1015), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1170), .B(KEYINPUT62), .C1(new_n1013), .C2(new_n1011), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1167), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1166), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n997), .B1(new_n1144), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n983), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  OR3_X1    g754(.A1(new_n1178), .A2(new_n1179), .A3(G1996), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n983), .B1(new_n986), .B2(new_n731), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1178), .B2(G1996), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT47), .Z(new_n1184));
  XOR2_X1   g759(.A(new_n989), .B(KEYINPUT125), .Z(new_n1185));
  NAND2_X1  g760(.A1(new_n988), .A2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n720), .A2(G2067), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1178), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n994), .A2(new_n983), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT48), .Z(new_n1190));
  AOI21_X1  g765(.A(new_n1190), .B1(new_n983), .B2(new_n991), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1184), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1177), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(G227), .A2(new_n460), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n669), .A2(new_n704), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1198), .A2(new_n970), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n882), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1200));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1200), .ZN(G308));
  INV_X1    g775(.A(G308), .ZN(G225));
endmodule


