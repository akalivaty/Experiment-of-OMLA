//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n203));
  INV_X1    g002(.A(G226gat), .ZN(new_n204));
  INV_X1    g003(.A(G233gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT23), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  AND4_X1   g011(.A1(KEYINPUT25), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(G190gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n218), .A2(new_n217), .B1(new_n214), .B2(G190gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT26), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n218), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT28), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT27), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT27), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G183gat), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT28), .A4(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n235), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n206), .B1(new_n228), .B2(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n219), .A2(new_n220), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n249), .A2(new_n224), .B1(new_n222), .B2(new_n213), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n240), .A2(new_n242), .A3(new_n237), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT28), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n243), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n235), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n250), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n204), .A2(new_n205), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n246), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G211gat), .ZN(new_n261));
  INV_X1    g060(.A(G218gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n263), .A2(KEYINPUT22), .ZN(new_n264));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(KEYINPUT22), .B2(new_n263), .ZN(new_n268));
  INV_X1    g067(.A(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n260), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n218), .B(new_n233), .C1(new_n230), .C2(new_n231), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT65), .B(new_n274), .C1(new_n254), .C2(new_n243), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n256), .B1(new_n255), .B2(new_n235), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n259), .B(new_n228), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n228), .A2(new_n245), .ZN(new_n278));
  INV_X1    g077(.A(new_n206), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n271), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n228), .A2(new_n259), .A3(new_n245), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n272), .B(new_n284), .C1(new_n258), .C2(new_n206), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n228), .B1(new_n275), .B2(new_n276), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n279), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n272), .A4(new_n284), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G8gat), .B(G36gat), .Z(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT73), .ZN(new_n293));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND3_X1  g094(.A1(new_n283), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT30), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n273), .A2(new_n282), .B1(new_n286), .B2(new_n290), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n295), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n286), .A2(new_n290), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT71), .B1(new_n281), .B2(new_n271), .ZN(new_n303));
  AOI211_X1 g102(.A(new_n202), .B(new_n272), .C1(new_n277), .C2(new_n280), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT72), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n283), .A2(new_n307), .A3(new_n291), .ZN(new_n308));
  INV_X1    g107(.A(new_n295), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G127gat), .A2(G134gat), .ZN(new_n312));
  INV_X1    g111(.A(G127gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT66), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G127gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n317), .B2(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G113gat), .B2(G120gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n312), .ZN(new_n325));
  NAND2_X1  g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n322), .A2(KEYINPUT67), .ZN(new_n329));
  OAI21_X1  g128(.A(G120gat), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n318), .A2(new_n324), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n333));
  AND2_X1   g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT74), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G141gat), .ZN(new_n337));
  INV_X1    g136(.A(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G155gat), .B(G162gat), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348));
  INV_X1    g147(.A(G155gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n346), .A2(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n339), .A2(KEYINPUT76), .A3(new_n341), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n331), .A2(new_n332), .A3(new_n345), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT80), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n318), .A2(new_n324), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n327), .A2(new_n330), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT4), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n343), .A2(new_n344), .B1(new_n353), .B2(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n332), .A4(new_n331), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n357), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT77), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n369), .A3(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n367), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n368), .A2(new_n370), .A3(new_n361), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n373), .B(KEYINPUT78), .Z(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT5), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n366), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n362), .B2(new_n356), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n372), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n363), .B(new_n331), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n374), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n378), .B2(new_n381), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n376), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(new_n389), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392));
  INV_X1    g191(.A(new_n389), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n376), .C1(new_n383), .C2(new_n384), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n311), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n287), .A2(new_n331), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n361), .B(new_n228), .C1(new_n275), .C2(new_n276), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT32), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G15gat), .B(G43gat), .Z(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n407), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n401), .B(KEYINPUT32), .C1(new_n403), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n400), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(new_n398), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT34), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(KEYINPUT68), .ZN(new_n416));
  AOI211_X1 g215(.A(new_n399), .B(new_n416), .C1(new_n397), .C2(new_n400), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n408), .A3(new_n410), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT31), .B(G50gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(G228gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n205), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT3), .B1(new_n271), .B2(new_n203), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n363), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n271), .B1(new_n371), .B2(new_n203), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n264), .A2(KEYINPUT81), .A3(new_n265), .A4(new_n266), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n203), .B(new_n433), .C1(new_n271), .C2(KEYINPUT81), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n363), .B1(new_n434), .B2(new_n367), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n435), .A2(new_n430), .B1(new_n426), .B2(new_n205), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n425), .B1(new_n437), .B2(G22gat), .ZN(new_n438));
  XOR2_X1   g237(.A(KEYINPUT82), .B(G22gat), .Z(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n432), .A2(new_n436), .A3(new_n442), .A4(new_n439), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n445));
  INV_X1    g244(.A(new_n439), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n434), .A2(new_n367), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n358), .ZN(new_n448));
  INV_X1    g247(.A(new_n430), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n427), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n450), .B2(new_n431), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n440), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n445), .B1(new_n452), .B2(new_n425), .ZN(new_n453));
  INV_X1    g252(.A(new_n425), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT83), .B(new_n454), .C1(new_n451), .C2(new_n440), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n444), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n396), .A2(new_n422), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT69), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n420), .A2(new_n458), .A3(new_n421), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n418), .A2(new_n408), .A3(KEYINPUT69), .A4(new_n410), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT35), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n461), .A2(new_n462), .A3(new_n456), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n457), .A2(KEYINPUT35), .B1(new_n463), .B2(new_n396), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n459), .A2(new_n466), .A3(new_n460), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n420), .A2(KEYINPUT36), .A3(new_n421), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n396), .B2(new_n456), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n380), .A2(new_n374), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n366), .A2(new_n372), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n374), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n474), .B(new_n476), .C1(new_n473), .C2(new_n472), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n471), .A3(new_n374), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n478), .A2(KEYINPUT86), .A3(new_n393), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT86), .B1(new_n478), .B2(new_n393), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT40), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n311), .A2(new_n391), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n485), .A2(new_n456), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n395), .A2(new_n390), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n295), .B1(new_n298), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n288), .A2(new_n284), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n490), .B2(new_n271), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n281), .A2(new_n272), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT38), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n489), .A2(new_n493), .B1(new_n298), .B2(new_n295), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT38), .ZN(new_n495));
  INV_X1    g294(.A(new_n489), .ZN(new_n496));
  INV_X1    g295(.A(new_n308), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n307), .B1(new_n283), .B2(new_n291), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n499), .B2(KEYINPUT37), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n487), .B(new_n494), .C1(new_n495), .C2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n465), .A2(new_n470), .B1(new_n486), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n469), .B(KEYINPUT85), .C1(new_n396), .C2(new_n456), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n464), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  NOR3_X1   g304(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT90), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n506), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n508), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n512), .B1(new_n520), .B2(new_n510), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n521), .B1(new_n516), .B2(new_n517), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n523), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n505), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT92), .B1(new_n532), .B2(new_n531), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n538), .B(KEYINPUT13), .Z(new_n543));
  NAND3_X1  g342(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n535), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n536), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n540), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G169gat), .B(G197gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT89), .ZN(new_n549));
  XOR2_X1   g348(.A(G113gat), .B(G141gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n540), .A2(new_n545), .A3(new_n554), .A4(new_n546), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n504), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n561));
  AND2_X1   g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n563));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567));
  INV_X1    g366(.A(new_n533), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  INV_X1    g371(.A(G92gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT96), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n570), .A2(new_n579), .A3(new_n576), .A4(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n532), .B2(KEYINPUT17), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n525), .A2(KEYINPUT97), .A3(new_n533), .A4(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT98), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n523), .A2(new_n581), .B1(KEYINPUT41), .B2(new_n562), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n586), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n566), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n565), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT9), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  INV_X1    g401(.A(G64gat), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n603), .A2(G57gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n604), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT9), .ZN(new_n612));
  NAND2_X1  g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT93), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(G71gat), .B2(G78gat), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n531), .B1(new_n619), .B2(new_n618), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT95), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n624), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n561), .B1(new_n598), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n581), .A2(new_n618), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n577), .A2(new_n618), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n610), .A4(new_n617), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G230gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n205), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n637), .A2(new_n645), .A3(new_n638), .ZN(new_n648));
  XOR2_X1   g447(.A(G120gat), .B(G148gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT100), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n645), .B1(new_n641), .B2(new_n642), .ZN(new_n655));
  INV_X1    g454(.A(new_n648), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n560), .A2(new_n635), .A3(new_n636), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n395), .A2(new_n390), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT101), .B(G1gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  AND2_X1   g463(.A1(new_n301), .A2(new_n310), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n530), .B2(new_n666), .ZN(new_n669));
  MUX2_X1   g468(.A(new_n668), .B(new_n669), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n660), .B2(new_n469), .ZN(new_n671));
  INV_X1    g470(.A(new_n461), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n660), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n660), .A2(new_n456), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NOR3_X1   g476(.A1(new_n597), .A2(new_n633), .A3(new_n658), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n560), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(G29gat), .A3(new_n661), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n682), .B(KEYINPUT44), .C1(new_n504), .C2(new_n597), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n467), .A2(new_n468), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n456), .B1(new_n661), .B2(new_n665), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n465), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n495), .B1(new_n687), .B2(new_n489), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n494), .A2(new_n395), .A3(new_n390), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n485), .B(new_n456), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n503), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n463), .A2(new_n396), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n661), .A2(new_n665), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n456), .A2(new_n421), .A3(new_n420), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT35), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n597), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT103), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT104), .B1(new_n396), .B2(new_n456), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n690), .A2(new_n700), .A3(new_n702), .A4(new_n469), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n597), .B1(new_n703), .B2(new_n696), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n698), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n633), .B(KEYINPUT102), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n558), .A2(new_n659), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n487), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G29gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n681), .A2(new_n712), .ZN(G1328gat));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n311), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G36gat), .ZN(new_n715));
  AOI211_X1 g514(.A(G36gat), .B(new_n665), .C1(KEYINPUT105), .C2(KEYINPUT46), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n560), .A2(new_n678), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n684), .A3(new_n709), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n679), .A2(G43gat), .A3(new_n672), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n721), .B(KEYINPUT47), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n722), .B2(G43gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(KEYINPUT106), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n725), .A2(new_n728), .ZN(G1330gat));
  INV_X1    g528(.A(new_n444), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n452), .A2(new_n425), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT83), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n452), .A2(new_n445), .A3(new_n425), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n706), .A2(new_n734), .A3(new_n709), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(new_n735), .B2(G50gat), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n679), .A2(G50gat), .A3(new_n456), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n735), .B2(G50gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI221_X4 g539(.A(new_n737), .B1(KEYINPUT107), .B2(KEYINPUT48), .C1(new_n735), .C2(G50gat), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n635), .A2(new_n636), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n743), .A2(new_n558), .A3(new_n659), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n703), .A2(new_n696), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n487), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g550(.A1(new_n747), .A2(new_n748), .A3(new_n665), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  AND2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n752), .B2(new_n753), .ZN(G1333gat));
  NAND3_X1  g555(.A1(new_n749), .A2(new_n599), .A3(new_n461), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n747), .A2(new_n748), .A3(new_n469), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n599), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n749), .A2(new_n734), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n558), .A2(new_n633), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n704), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT109), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n572), .A3(new_n487), .A4(new_n658), .ZN(new_n771));
  INV_X1    g570(.A(new_n764), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n659), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n706), .A2(new_n487), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n572), .B2(new_n774), .ZN(G1336gat));
  NOR3_X1   g574(.A1(new_n659), .A2(new_n665), .A3(G92gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n706), .A2(new_n311), .A3(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT110), .B1(new_n778), .B2(G92gat), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n597), .B(new_n772), .C1(new_n703), .C2(new_n696), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n766), .B1(new_n784), .B2(KEYINPUT111), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n765), .A2(new_n786), .A3(KEYINPUT51), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n787), .A3(new_n776), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT112), .A4(new_n776), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n782), .A2(new_n783), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n781), .B1(new_n793), .B2(new_n780), .ZN(G1337gat));
  NOR3_X1   g593(.A1(new_n672), .A2(G99gat), .A3(new_n659), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n706), .A2(new_n684), .A3(new_n773), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G99gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1338gat));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n659), .A2(new_n456), .A3(G106gat), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n770), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n800), .B1(new_n770), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n706), .A2(new_n734), .A3(new_n773), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n785), .A2(new_n787), .A3(new_n802), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n805), .A2(new_n809), .B1(new_n811), .B2(new_n808), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n641), .A2(new_n645), .A3(new_n642), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n653), .B1(new_n655), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n654), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n815), .B2(new_n817), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n820), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(KEYINPUT115), .A3(new_n654), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n823), .A3(new_n558), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n537), .B2(new_n539), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n826), .B(new_n538), .C1(new_n534), .C2(new_n536), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n557), .B(new_n658), .C1(new_n829), .C2(new_n553), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n598), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n821), .A2(new_n823), .ZN(new_n832));
  INV_X1    g631(.A(new_n553), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n825), .A2(new_n828), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n827), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n557), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n832), .A2(new_n836), .A3(new_n597), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n707), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n635), .A2(new_n559), .A3(new_n636), .A4(new_n659), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n734), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n661), .A2(new_n311), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n461), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n559), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n661), .B1(new_n838), .B2(new_n839), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n694), .A2(new_n311), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n328), .A2(new_n329), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n558), .A2(new_n855), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n845), .A2(new_n846), .B1(new_n854), .B2(new_n856), .ZN(G1340gat));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n658), .A2(new_n323), .ZN(new_n859));
  INV_X1    g658(.A(new_n853), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n851), .ZN(new_n861));
  OAI21_X1  g660(.A(G120gat), .B1(new_n842), .B2(new_n659), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT119), .B(new_n862), .C1(new_n854), .C2(new_n859), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(new_n317), .B1(new_n842), .B2(new_n707), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n633), .A2(new_n314), .A3(new_n316), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n849), .B2(new_n868), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n597), .A2(G134gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n847), .A2(new_n848), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n842), .B2(new_n597), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT120), .ZN(G1343gat));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n835), .A2(new_n878), .A3(new_n557), .A4(new_n658), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n830), .A2(KEYINPUT121), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n819), .A2(new_n820), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n558), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n836), .A2(new_n597), .ZN(new_n884));
  INV_X1    g683(.A(new_n832), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n883), .A2(new_n597), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n839), .B1(new_n886), .B2(new_n633), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n877), .B1(new_n887), .B2(new_n734), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT57), .B(new_n456), .C1(new_n838), .C2(new_n839), .ZN(new_n889));
  INV_X1    g688(.A(new_n841), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n684), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n559), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n684), .A2(new_n311), .A3(new_n456), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n847), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(G141gat), .A3(new_n559), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n337), .B1(new_n901), .B2(new_n558), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT58), .B1(new_n902), .B2(new_n898), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1344gat));
  INV_X1    g703(.A(new_n897), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n338), .A3(new_n658), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n338), .C1(new_n901), .C2(new_n658), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n838), .A2(new_n839), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n734), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n743), .A2(new_n558), .A3(new_n658), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n883), .A2(new_n597), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n884), .A2(new_n881), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n633), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n877), .B(new_n734), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n911), .A2(new_n658), .A3(new_n891), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n908), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n906), .B1(new_n907), .B2(new_n918), .ZN(G1345gat));
  NOR3_X1   g718(.A1(new_n893), .A2(new_n349), .A3(new_n707), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n897), .B2(new_n634), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n897), .A2(KEYINPUT122), .A3(new_n634), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(G155gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n893), .B2(new_n597), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n350), .A3(new_n598), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n487), .A2(new_n665), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n461), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n840), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n207), .A3(new_n559), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT123), .B1(new_n909), .B2(new_n661), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n934), .B(new_n487), .C1(new_n838), .C2(new_n839), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n694), .A2(new_n665), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n558), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n932), .B1(new_n938), .B2(new_n207), .ZN(G1348gat));
  OAI21_X1  g738(.A(G176gat), .B1(new_n931), .B2(new_n659), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n658), .A2(new_n208), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1349gat));
  NAND2_X1  g742(.A1(new_n633), .A2(new_n236), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n937), .B(new_n945), .C1(new_n933), .C2(new_n935), .ZN(new_n946));
  OAI21_X1  g745(.A(G183gat), .B1(new_n931), .B2(new_n707), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g748(.A1(new_n597), .A2(G190gat), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n937), .B(new_n950), .C1(new_n933), .C2(new_n935), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n840), .A2(new_n598), .A3(new_n930), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(G190gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n952), .B2(G190gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT125), .ZN(G1351gat));
  AND2_X1   g756(.A1(new_n928), .A2(new_n469), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n911), .A2(new_n916), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n559), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n684), .A2(new_n665), .A3(new_n456), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n936), .A2(KEYINPUT126), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n933), .B2(new_n935), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n558), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n961), .B1(new_n967), .B2(new_n960), .ZN(G1352gat));
  OR2_X1    g767(.A1(new_n659), .A2(G204gat), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT62), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT127), .B1(new_n959), .B2(new_n659), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G204gat), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n959), .A2(KEYINPUT127), .A3(new_n659), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n970), .B(new_n971), .C1(new_n973), .C2(new_n974), .ZN(G1353gat));
  NAND4_X1  g774(.A1(new_n963), .A2(new_n261), .A3(new_n633), .A4(new_n966), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n911), .A2(new_n633), .A3(new_n916), .A4(new_n958), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  NAND4_X1  g780(.A1(new_n963), .A2(new_n262), .A3(new_n598), .A4(new_n966), .ZN(new_n982));
  OAI21_X1  g781(.A(G218gat), .B1(new_n959), .B2(new_n597), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


