//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949;
  OR2_X1    g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT64), .B1(new_n189), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n188), .A3(new_n187), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT0), .A3(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(KEYINPUT64), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n202), .A3(G128), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n190), .A3(G143), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n192), .B(G146), .C1(new_n204), .C2(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G224), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G953), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n211), .B(new_n215), .C1(KEYINPUT85), .C2(new_n213), .ZN(new_n216));
  XOR2_X1   g030(.A(G110), .B(G122), .Z(new_n217));
  XOR2_X1   g031(.A(new_n217), .B(KEYINPUT8), .Z(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n219), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G116), .B(G119), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n220), .A3(new_n221), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT78), .B(G101), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n230), .B2(G107), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n229), .A2(new_n231), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n231), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n230), .A2(G107), .ZN(new_n238));
  OAI21_X1  g052(.A(G101), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n226), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n228), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n225), .B(KEYINPUT84), .Z(new_n245));
  NAND2_X1  g059(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n245), .A2(new_n246), .B1(new_n226), .B2(new_n242), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n218), .B(new_n244), .C1(new_n247), .C2(new_n240), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n235), .A2(new_n234), .A3(new_n231), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n236), .ZN(new_n251));
  INV_X1    g065(.A(new_n226), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n241), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n243), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n255), .A3(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n228), .A2(new_n236), .A3(new_n243), .A4(new_n239), .ZN(new_n258));
  INV_X1    g072(.A(new_n217), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT7), .B(new_n214), .C1(new_n210), .C2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n216), .A2(new_n248), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n210), .B(new_n214), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n257), .A2(KEYINPUT81), .A3(new_n258), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT81), .B1(new_n257), .B2(new_n258), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n217), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n260), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n257), .A2(new_n258), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT81), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n259), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT82), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n276), .B(new_n217), .C1(new_n267), .C2(new_n268), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n266), .B(new_n270), .C1(new_n277), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT83), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n276), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n279), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT83), .A3(new_n266), .A4(new_n270), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n265), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT86), .Z(new_n290));
  XOR2_X1   g104(.A(new_n290), .B(KEYINPUT87), .Z(new_n291));
  NOR2_X1   g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n290), .B(new_n265), .C1(new_n283), .C2(new_n287), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n296));
  INV_X1    g110(.A(new_n195), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n196), .B2(new_n198), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n300), .A2(KEYINPUT67), .A3(new_n195), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n251), .B(new_n256), .C1(new_n298), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT11), .ZN(new_n303));
  INV_X1    g117(.A(G134), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(G137), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(G137), .ZN(new_n306));
  INV_X1    g120(.A(G137), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT11), .A3(G134), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G131), .ZN(new_n310));
  INV_X1    g124(.A(G131), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n305), .A2(new_n308), .A3(new_n311), .A4(new_n306), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n207), .A2(new_n236), .A3(new_n239), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n316), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n302), .A2(new_n314), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n240), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n314), .B1(new_n322), .B2(new_n315), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT12), .B1(new_n313), .B2(KEYINPUT79), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G140), .ZN(new_n326));
  INV_X1    g140(.A(G227), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(G953), .ZN(new_n328));
  XOR2_X1   g142(.A(new_n326), .B(new_n328), .Z(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n320), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n302), .A2(new_n317), .A3(new_n318), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n313), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n333), .B2(new_n319), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G469), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n264), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n330), .B1(new_n320), .B2(new_n325), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n319), .A3(new_n329), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(G469), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(G469), .A2(G902), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G221), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT9), .B(G234), .Z(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(new_n264), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G214), .B1(G237), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n294), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G234), .ZN(new_n351));
  OAI21_X1  g165(.A(G217), .B1(new_n351), .B2(G902), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT72), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT22), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(new_n307), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n204), .A2(G119), .B1(KEYINPUT74), .B2(KEYINPUT23), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n204), .A2(G119), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G110), .ZN(new_n364));
  INV_X1    g178(.A(G119), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G128), .ZN(new_n366));
  AND2_X1   g180(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n367));
  NOR2_X1   g181(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n363), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT24), .B(G110), .Z(new_n371));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n366), .B2(new_n362), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n204), .A2(G119), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n365), .A2(G128), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT73), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n360), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n208), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G125), .A2(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT16), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(G146), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT24), .B(G110), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT73), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT73), .B1(new_n374), .B2(new_n375), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n363), .A2(new_n364), .A3(new_n369), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(KEYINPUT76), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n382), .A2(new_n190), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n378), .A2(new_n386), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT77), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n380), .B2(new_n381), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n397), .A2(new_n190), .A3(new_n384), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(new_n391), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n360), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n400), .A2(new_n401), .A3(new_n392), .A4(new_n393), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n190), .B1(new_n397), .B2(new_n384), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT75), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n386), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT75), .B(new_n190), .C1(new_n397), .C2(new_n384), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n363), .A2(new_n369), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G110), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n373), .A2(new_n376), .A3(new_n371), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n406), .A2(new_n407), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n359), .B1(new_n403), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n411), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n413), .B(new_n358), .C1(new_n395), .C2(new_n402), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT25), .B1(new_n415), .B2(new_n264), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n417));
  NOR4_X1   g231(.A1(new_n412), .A2(new_n414), .A3(new_n417), .A4(G902), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n354), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n394), .A2(KEYINPUT77), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n392), .A2(new_n393), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n401), .B1(new_n421), .B2(new_n400), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n411), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n358), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n403), .A2(new_n411), .A3(new_n359), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n264), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n419), .B1(new_n354), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n307), .A2(G134), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n304), .A2(G137), .ZN(new_n429));
  OAI21_X1  g243(.A(G131), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n312), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n207), .B1(new_n313), .B2(new_n200), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT66), .B1(new_n434), .B2(KEYINPUT30), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n313), .B1(new_n298), .B2(new_n301), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT68), .B1(new_n321), .B2(new_n431), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n312), .A2(new_n430), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n207), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT30), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n432), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n431), .A2(KEYINPUT65), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n207), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n200), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(new_n314), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n435), .A2(new_n442), .A3(new_n254), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n254), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n436), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(G101), .ZN(new_n455));
  NOR2_X1   g269(.A1(G237), .A2(G953), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G210), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n451), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT31), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n451), .A2(KEYINPUT31), .A3(new_n453), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n200), .A2(new_n295), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT67), .B1(new_n300), .B2(new_n195), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n314), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n321), .A2(new_n431), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n466), .A2(new_n254), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT28), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n447), .A2(new_n254), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n453), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n458), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT32), .ZN(new_n477));
  INV_X1    g291(.A(G472), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n264), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n461), .A2(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n264), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT32), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n451), .A2(new_n453), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n474), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(KEYINPUT70), .A3(new_n474), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n437), .A2(new_n440), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n254), .B1(new_n466), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n453), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT71), .A4(new_n452), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n469), .B1(new_n497), .B2(KEYINPUT28), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n474), .A2(new_n488), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G472), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n427), .B1(new_n483), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n456), .A2(G143), .A3(G214), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G143), .B1(new_n456), .B2(G214), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n456), .A2(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n192), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n311), .A3(new_n504), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n398), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n382), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n513));
  OR2_X1    g327(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n382), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n190), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n505), .A2(new_n506), .ZN(new_n519));
  NAND2_X1  g333(.A1(KEYINPUT18), .A2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n512), .A2(G146), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n393), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n311), .B1(new_n509), .B2(new_n504), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT18), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n511), .A2(new_n518), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G113), .B(G122), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n230), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT89), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n406), .A2(new_n407), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n507), .A2(new_n531), .A3(new_n510), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n519), .A2(new_n520), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n393), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n524), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n527), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n510), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n386), .B1(new_n538), .B2(new_n523), .ZN(new_n539));
  AOI21_X1  g353(.A(G146), .B1(new_n515), .B2(new_n516), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n542));
  INV_X1    g356(.A(new_n527), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n528), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G475), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n264), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT20), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n547), .A2(KEYINPUT20), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT91), .B(G475), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n533), .A2(new_n536), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n527), .A2(KEYINPUT92), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n557), .B2(G902), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(G234), .A2(G237), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(G952), .A3(new_n355), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT21), .B(G898), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(G902), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT94), .B(KEYINPUT15), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT95), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OR3_X1    g387(.A1(new_n571), .A2(KEYINPUT95), .A3(new_n572), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n573), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n344), .A2(G217), .A3(new_n355), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G122), .ZN(new_n578));
  OR3_X1    g392(.A1(new_n578), .A2(KEYINPUT93), .A3(G116), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT93), .B1(new_n578), .B2(G116), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n579), .A2(new_n580), .B1(G116), .B2(new_n578), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(G116), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n233), .B1(new_n582), .B2(KEYINPUT14), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G128), .B(G143), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n304), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(KEYINPUT13), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n204), .A2(KEYINPUT13), .A3(G143), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n304), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n588), .A2(new_n590), .B1(new_n304), .B2(new_n585), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n581), .A2(new_n233), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n581), .A2(new_n233), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n577), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n587), .A2(new_n594), .A3(new_n577), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  MUX2_X1   g412(.A(new_n573), .B(new_n575), .S(new_n598), .Z(new_n599));
  NOR2_X1   g413(.A1(new_n570), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n350), .A2(new_n503), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n601), .B(new_n229), .Z(G3));
  INV_X1    g416(.A(new_n290), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n283), .A2(new_n287), .ZN(new_n604));
  INV_X1    g418(.A(new_n265), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n348), .B1(new_n606), .B2(new_n293), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT97), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n348), .C1(new_n606), .C2(new_n293), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n568), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n598), .A2(new_n572), .ZN(new_n614));
  NAND2_X1  g428(.A1(G478), .A2(G902), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n597), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n597), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n595), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n596), .B(new_n597), .C1(new_n617), .C2(new_n616), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n614), .B(new_n615), .C1(new_n622), .C2(new_n572), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n560), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n476), .A2(new_n478), .A3(new_n264), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n480), .B2(G902), .ZN(new_n627));
  INV_X1    g441(.A(new_n427), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n347), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT96), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(new_n552), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n549), .A2(new_n551), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n637), .B2(new_n636), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(new_n558), .A3(new_n599), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n613), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n631), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n233), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G9));
  INV_X1    g459(.A(new_n600), .ZN(new_n646));
  INV_X1    g460(.A(new_n347), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n288), .A2(new_n603), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n291), .B2(new_n288), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n348), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n626), .A2(new_n627), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n426), .A2(new_n417), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n424), .A2(KEYINPUT25), .A3(new_n264), .A4(new_n425), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n353), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n423), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n264), .A3(new_n353), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n419), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n646), .A2(new_n650), .A3(new_n651), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT102), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT37), .B(G110), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n662), .B1(new_n483), .B2(new_n502), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n647), .A3(new_n610), .A4(new_n608), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT103), .B(G900), .Z(new_n670));
  AOI21_X1  g484(.A(new_n563), .B1(new_n670), .B2(new_n567), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n639), .A2(new_n558), .A3(new_n599), .A4(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n667), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n479), .A2(new_n482), .B1(new_n501), .B2(G472), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n675), .A2(new_n347), .A3(new_n662), .ZN(new_n676));
  INV_X1    g490(.A(new_n673), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n611), .A2(new_n676), .A3(new_n677), .A4(KEYINPUT104), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  NAND2_X1  g494(.A1(new_n497), .A2(new_n474), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n459), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n264), .B1(new_n682), .B2(KEYINPUT105), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(KEYINPUT105), .B2(new_n682), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(new_n478), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n483), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n348), .A3(new_n662), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n671), .B(KEYINPUT39), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n647), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n687), .B1(KEYINPUT40), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n294), .B(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n694));
  INV_X1    g508(.A(new_n599), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n560), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n693), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  NAND2_X1  g512(.A1(new_n668), .A2(new_n647), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n560), .A2(new_n623), .A3(new_n671), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n608), .A2(new_n700), .A3(new_n610), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n699), .B1(new_n701), .B2(KEYINPUT106), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n611), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NAND2_X1  g520(.A1(new_n335), .A2(new_n264), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n346), .A3(new_n337), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n675), .A2(new_n427), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n613), .A2(new_n624), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND4_X1  g527(.A1(new_n611), .A2(new_n710), .A3(new_n640), .A4(new_n569), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NOR2_X1   g529(.A1(new_n612), .A2(new_n709), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n600), .A3(new_n668), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  OAI21_X1  g532(.A(new_n463), .B1(new_n498), .B2(new_n458), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n478), .A3(new_n264), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n627), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n628), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n568), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n716), .A2(new_n696), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  INV_X1    g539(.A(new_n709), .ZN(new_n726));
  INV_X1    g540(.A(new_n662), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n611), .A2(new_n700), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NOR2_X1   g544(.A1(new_n649), .A2(new_n349), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n503), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n341), .B(KEYINPUT107), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n340), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n345), .B1(new_n337), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n624), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n732), .A2(new_n740), .A3(new_n733), .A4(new_n737), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n737), .A2(new_n503), .A3(new_n672), .A4(new_n731), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n739), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND3_X1  g560(.A1(new_n732), .A2(new_n677), .A3(new_n736), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NAND2_X1  g562(.A1(new_n338), .A2(new_n339), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G469), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n734), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n734), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n337), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n346), .A3(new_n689), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n559), .A2(new_n623), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n651), .A4(new_n727), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n765), .B(new_n731), .C1(new_n764), .C2(new_n763), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT111), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  NAND2_X1  g582(.A1(new_n756), .A2(new_n346), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT47), .Z(new_n770));
  NAND2_X1  g584(.A1(new_n731), .A2(new_n672), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n624), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n675), .A2(new_n427), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT112), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  OR2_X1    g591(.A1(new_n760), .A2(new_n562), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n649), .A2(new_n709), .A3(new_n349), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n503), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT48), .Z(new_n782));
  NOR2_X1   g596(.A1(new_n778), .A2(new_n722), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n349), .A3(new_n692), .A4(new_n726), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT50), .Z(new_n785));
  NAND3_X1  g599(.A1(new_n779), .A2(new_n728), .A3(new_n780), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n708), .A2(new_n337), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n346), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n731), .B(new_n783), .C1(new_n770), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n686), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n780), .A3(new_n628), .A4(new_n563), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n560), .A2(new_n623), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n785), .A2(new_n786), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  AND4_X1   g611(.A1(G952), .A2(new_n796), .A3(new_n355), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n624), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n568), .B(new_n623), .C1(new_n553), .C2(new_n558), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n649), .A2(new_n348), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n649), .A2(KEYINPUT113), .A3(new_n348), .A4(new_n801), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n630), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n601), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n714), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n601), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n663), .B1(new_n810), .B2(KEYINPUT114), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n811), .A3(new_n717), .A4(new_n724), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n745), .A2(new_n747), .ZN(new_n813));
  OR4_X1    g627(.A1(new_n570), .A2(new_n650), .A3(new_n695), .A4(new_n629), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n711), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n676), .A2(new_n558), .A3(new_n695), .A4(new_n639), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n728), .A2(new_n737), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n771), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n608), .A2(new_n610), .A3(new_n696), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n736), .A2(new_n419), .A3(new_n657), .A4(new_n672), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n820), .A2(new_n686), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n679), .A2(new_n705), .A3(new_n729), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n674), .A2(new_n678), .B1(new_n702), .B2(new_n704), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n729), .A4(new_n825), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n819), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n832), .A2(KEYINPUT53), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT54), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n838), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n831), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n798), .A2(new_n800), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n782), .B(new_n845), .C1(new_n716), .C2(new_n783), .ZN(new_n846));
  NOR2_X1   g660(.A1(G952), .A2(G953), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n790), .A2(new_n628), .A3(new_n348), .A4(new_n758), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n787), .B(KEYINPUT49), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n692), .A2(new_n849), .A3(new_n346), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n846), .A2(new_n847), .B1(new_n848), .B2(new_n850), .ZN(G75));
  NAND2_X1  g665(.A1(new_n286), .A2(new_n270), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(new_n266), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT55), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n828), .A2(new_n834), .A3(new_n830), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n834), .B1(new_n828), .B2(new_n830), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n837), .B1(new_n857), .B2(new_n819), .ZN(new_n858));
  INV_X1    g672(.A(new_n843), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n264), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n290), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT56), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n854), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n355), .A2(G952), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n854), .A2(new_n863), .ZN(new_n866));
  INV_X1    g680(.A(new_n291), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(G51));
  OAI21_X1  g683(.A(KEYINPUT54), .B1(new_n858), .B2(new_n859), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(new_n844), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n860), .A2(KEYINPUT119), .A3(new_n842), .ZN(new_n873));
  XNOR2_X1  g687(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n734), .B(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n876), .A2(KEYINPUT120), .A3(new_n335), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT120), .B1(new_n876), .B2(new_n335), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n861), .A2(G469), .A3(new_n750), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n865), .B1(new_n879), .B2(new_n880), .ZN(G54));
  NAND2_X1  g695(.A1(new_n841), .A2(new_n843), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n883));
  INV_X1    g697(.A(new_n545), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n865), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT121), .ZN(G60));
  XOR2_X1   g703(.A(new_n615), .B(KEYINPUT59), .Z(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n840), .B2(new_n844), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n886), .B1(new_n891), .B2(new_n622), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n620), .B2(new_n621), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n872), .A2(new_n873), .A3(new_n893), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT122), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n892), .B2(new_n894), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(G63));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT124), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT60), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n860), .A2(new_n900), .B1(new_n414), .B2(new_n412), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n860), .A2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(new_n656), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n886), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g721(.A(new_n812), .ZN(new_n908));
  INV_X1    g722(.A(new_n815), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n355), .ZN(new_n911));
  OAI21_X1  g725(.A(G953), .B1(new_n565), .B2(new_n212), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT125), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n852), .B1(G898), .B2(new_n355), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G69));
  AND2_X1   g730(.A1(new_n745), .A2(new_n747), .ZN(new_n917));
  INV_X1    g731(.A(new_n757), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n503), .A3(new_n820), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n766), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n829), .A2(new_n729), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n773), .B2(new_n774), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT126), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n355), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n435), .A2(new_n442), .A3(new_n450), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(new_n517), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n327), .A2(G900), .A3(G953), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n930));
  INV_X1    g744(.A(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n921), .A2(new_n697), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n775), .B1(KEYINPUT62), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n624), .B1(new_n560), .B2(new_n599), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n690), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n732), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n933), .A2(new_n934), .A3(new_n766), .A4(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n930), .B(new_n931), .C1(new_n938), .C2(G953), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n939), .ZN(G72));
  NAND2_X1  g754(.A1(G472), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT63), .Z(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n924), .B2(new_n910), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(new_n453), .A3(new_n474), .A4(new_n451), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n938), .B2(new_n910), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n458), .A3(new_n484), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n487), .A2(new_n459), .A3(new_n490), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n839), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n944), .A2(new_n886), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT127), .ZN(G57));
endmodule


