

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578;

  XOR2_X1 U320 ( .A(n313), .B(n312), .Z(n288) );
  XNOR2_X1 U321 ( .A(KEYINPUT108), .B(KEYINPUT48), .ZN(n369) );
  XNOR2_X1 U322 ( .A(n370), .B(n369), .ZN(n515) );
  INV_X1 U323 ( .A(n373), .ZN(n319) );
  XNOR2_X1 U324 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U325 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U326 ( .A(KEYINPUT120), .B(n442), .ZN(n560) );
  XNOR2_X1 U327 ( .A(n444), .B(KEYINPUT58), .ZN(n445) );
  XNOR2_X1 U328 ( .A(n446), .B(n445), .ZN(G1351GAT) );
  XNOR2_X1 U329 ( .A(G36GAT), .B(G190GAT), .ZN(n289) );
  XNOR2_X1 U330 ( .A(n289), .B(KEYINPUT78), .ZN(n377) );
  XOR2_X1 U331 ( .A(n377), .B(KEYINPUT10), .Z(n291) );
  XOR2_X1 U332 ( .A(G50GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U333 ( .A(n415), .B(G218GAT), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n297) );
  XOR2_X1 U335 ( .A(G92GAT), .B(KEYINPUT75), .Z(n293) );
  XNOR2_X1 U336 ( .A(G99GAT), .B(G85GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n326) );
  XOR2_X1 U338 ( .A(n326), .B(G106GAT), .Z(n295) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n305) );
  XOR2_X1 U342 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n299) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U345 ( .A(KEYINPUT73), .B(n300), .Z(n343) );
  XOR2_X1 U346 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n302) );
  XNOR2_X1 U347 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n343), .B(n303), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n547) );
  INV_X1 U351 ( .A(n547), .ZN(n443) );
  XOR2_X1 U352 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n307) );
  XNOR2_X1 U353 ( .A(KEYINPUT83), .B(KEYINPUT14), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n324) );
  XOR2_X1 U355 ( .A(G155GAT), .B(G211GAT), .Z(n309) );
  XNOR2_X1 U356 ( .A(G127GAT), .B(G71GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U358 ( .A(KEYINPUT82), .B(G64GAT), .Z(n311) );
  XNOR2_X1 U359 ( .A(G22GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n315) );
  NAND2_X1 U362 ( .A1(G231GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U364 ( .A(KEYINPUT81), .B(n316), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n288), .B(n317), .ZN(n322) );
  XNOR2_X1 U366 ( .A(G15GAT), .B(G1GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n318), .B(KEYINPUT74), .ZN(n339) );
  XOR2_X1 U368 ( .A(G57GAT), .B(KEYINPUT13), .Z(n325) );
  XNOR2_X1 U369 ( .A(n339), .B(n325), .ZN(n320) );
  XOR2_X1 U370 ( .A(G8GAT), .B(G183GAT), .Z(n373) );
  XOR2_X1 U371 ( .A(n324), .B(n323), .Z(n571) );
  INV_X1 U372 ( .A(n571), .ZN(n543) );
  XNOR2_X1 U373 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n338) );
  XOR2_X1 U374 ( .A(n326), .B(n325), .Z(n330) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n419) );
  XOR2_X1 U378 ( .A(G176GAT), .B(G64GAT), .Z(n374) );
  XNOR2_X1 U379 ( .A(n419), .B(n374), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n337) );
  XOR2_X1 U381 ( .A(G120GAT), .B(G71GAT), .Z(n424) );
  XOR2_X1 U382 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n332) );
  XNOR2_X1 U383 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n424), .B(n333), .Z(n335) );
  NAND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n363) );
  XOR2_X1 U389 ( .A(n338), .B(n363), .Z(n557) );
  INV_X1 U390 ( .A(n557), .ZN(n538) );
  XOR2_X1 U391 ( .A(G141GAT), .B(G22GAT), .Z(n416) );
  XOR2_X1 U392 ( .A(n339), .B(n416), .Z(n341) );
  XNOR2_X1 U393 ( .A(G50GAT), .B(G36GAT), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n356) );
  XOR2_X1 U396 ( .A(KEYINPUT30), .B(G197GAT), .Z(n345) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G113GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U399 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n347) );
  XNOR2_X1 U400 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U402 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U403 ( .A(G8GAT), .B(KEYINPUT68), .Z(n351) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U406 ( .A(KEYINPUT71), .B(n352), .ZN(n353) );
  XOR2_X1 U407 ( .A(n354), .B(n353), .Z(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n564) );
  INV_X1 U409 ( .A(n564), .ZN(n535) );
  NAND2_X1 U410 ( .A1(n538), .A2(n535), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n357), .B(KEYINPUT46), .ZN(n358) );
  XNOR2_X1 U412 ( .A(KEYINPUT106), .B(n358), .ZN(n359) );
  NAND2_X1 U413 ( .A1(n359), .A2(n443), .ZN(n360) );
  NOR2_X1 U414 ( .A1(n543), .A2(n360), .ZN(n361) );
  XNOR2_X1 U415 ( .A(KEYINPUT47), .B(n361), .ZN(n368) );
  XOR2_X1 U416 ( .A(KEYINPUT36), .B(n547), .Z(n575) );
  NOR2_X1 U417 ( .A1(n571), .A2(n575), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n362), .B(KEYINPUT45), .ZN(n364) );
  NAND2_X1 U419 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n365), .B(KEYINPUT107), .ZN(n366) );
  NAND2_X1 U421 ( .A1(n366), .A2(n564), .ZN(n367) );
  NAND2_X1 U422 ( .A1(n368), .A2(n367), .ZN(n370) );
  XOR2_X1 U423 ( .A(G211GAT), .B(KEYINPUT21), .Z(n372) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(G218GAT), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n420) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n384) );
  XOR2_X1 U427 ( .A(G92GAT), .B(KEYINPUT91), .Z(n376) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U430 ( .A(n378), .B(n377), .Z(n382) );
  XOR2_X1 U431 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n380) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n425) );
  XNOR2_X1 U434 ( .A(n425), .B(G204GAT), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U437 ( .A(n420), .B(n385), .Z(n473) );
  AND2_X1 U438 ( .A1(n515), .A2(n473), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n386), .B(KEYINPUT54), .ZN(n406) );
  XOR2_X1 U440 ( .A(G127GAT), .B(KEYINPUT0), .Z(n388) );
  XNOR2_X1 U441 ( .A(G113GAT), .B(G134GAT), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n428) );
  XOR2_X1 U443 ( .A(KEYINPUT90), .B(n428), .Z(n390) );
  NAND2_X1 U444 ( .A1(G225GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n405) );
  XOR2_X1 U446 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U447 ( .A(G29GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U449 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n394) );
  XNOR2_X1 U450 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U452 ( .A(n396), .B(n395), .Z(n403) );
  XOR2_X1 U453 ( .A(G155GAT), .B(KEYINPUT2), .Z(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n408) );
  XOR2_X1 U456 ( .A(G57GAT), .B(G148GAT), .Z(n400) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(G1GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n408), .B(n401), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U461 ( .A(n405), .B(n404), .Z(n506) );
  NAND2_X1 U462 ( .A1(n406), .A2(n506), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n407), .B(KEYINPUT65), .ZN(n562) );
  XOR2_X1 U464 ( .A(KEYINPUT24), .B(n408), .Z(n410) );
  NAND2_X1 U465 ( .A1(G228GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n412) );
  XNOR2_X1 U468 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U473 ( .A(n420), .B(n419), .Z(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n458) );
  NAND2_X1 U475 ( .A1(n562), .A2(n458), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT55), .ZN(n441) );
  XOR2_X1 U477 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U478 ( .A(G43GAT), .B(G99GAT), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n432) );
  XOR2_X1 U480 ( .A(n428), .B(G176GAT), .Z(n430) );
  NAND2_X1 U481 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U483 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U484 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n434) );
  XNOR2_X1 U485 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U487 ( .A(KEYINPUT84), .B(G183GAT), .Z(n436) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(KEYINPUT66), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U491 ( .A(n440), .B(n439), .Z(n520) );
  INV_X1 U492 ( .A(n520), .ZN(n457) );
  NAND2_X1 U493 ( .A1(n441), .A2(n457), .ZN(n442) );
  NOR2_X1 U494 ( .A1(n443), .A2(n560), .ZN(n446) );
  INV_X1 U495 ( .A(G190GAT), .ZN(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n448) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n472) );
  NAND2_X1 U499 ( .A1(n535), .A2(n363), .ZN(n483) );
  NOR2_X1 U500 ( .A1(n571), .A2(n547), .ZN(n449) );
  XNOR2_X1 U501 ( .A(KEYINPUT16), .B(n449), .ZN(n469) );
  XOR2_X1 U502 ( .A(KEYINPUT27), .B(n473), .Z(n460) );
  NOR2_X1 U503 ( .A1(n506), .A2(n460), .ZN(n516) );
  XOR2_X1 U504 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n450) );
  XNOR2_X1 U505 ( .A(n458), .B(n450), .ZN(n518) );
  NAND2_X1 U506 ( .A1(n516), .A2(n518), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT92), .B(n451), .ZN(n452) );
  NOR2_X1 U508 ( .A1(n457), .A2(n452), .ZN(n453) );
  XNOR2_X1 U509 ( .A(KEYINPUT93), .B(n453), .ZN(n467) );
  NAND2_X1 U510 ( .A1(n473), .A2(n457), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n454), .A2(n458), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT25), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT95), .B(n456), .ZN(n464) );
  NOR2_X1 U514 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT26), .ZN(n563) );
  INV_X1 U516 ( .A(n460), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n563), .A2(n461), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT94), .B(n462), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n465), .A2(n506), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n468), .B(KEYINPUT96), .ZN(n480) );
  NAND2_X1 U523 ( .A1(n469), .A2(n480), .ZN(n494) );
  NOR2_X1 U524 ( .A1(n483), .A2(n494), .ZN(n470) );
  XNOR2_X1 U525 ( .A(KEYINPUT97), .B(n470), .ZN(n477) );
  NOR2_X1 U526 ( .A1(n506), .A2(n477), .ZN(n471) );
  XOR2_X1 U527 ( .A(n472), .B(n471), .Z(G1324GAT) );
  INV_X1 U528 ( .A(n473), .ZN(n509) );
  NOR2_X1 U529 ( .A1(n509), .A2(n477), .ZN(n474) );
  XOR2_X1 U530 ( .A(G8GAT), .B(n474), .Z(G1325GAT) );
  NOR2_X1 U531 ( .A1(n520), .A2(n477), .ZN(n476) );
  XNOR2_X1 U532 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  NOR2_X1 U534 ( .A1(n518), .A2(n477), .ZN(n478) );
  XOR2_X1 U535 ( .A(G22GAT), .B(n478), .Z(G1327GAT) );
  XOR2_X1 U536 ( .A(G29GAT), .B(KEYINPUT100), .Z(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT39), .B(n479), .ZN(n486) );
  NAND2_X1 U538 ( .A1(n571), .A2(n480), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n481), .A2(n575), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(KEYINPUT37), .ZN(n505) );
  NOR2_X1 U541 ( .A1(n505), .A2(n483), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT38), .B(n484), .Z(n492) );
  NOR2_X1 U543 ( .A1(n506), .A2(n492), .ZN(n485) );
  XOR2_X1 U544 ( .A(n486), .B(n485), .Z(G1328GAT) );
  NOR2_X1 U545 ( .A1(n492), .A2(n509), .ZN(n487) );
  XOR2_X1 U546 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n489) );
  XNOR2_X1 U548 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n491) );
  NOR2_X1 U550 ( .A1(n492), .A2(n520), .ZN(n490) );
  XOR2_X1 U551 ( .A(n491), .B(n490), .Z(G1330GAT) );
  NOR2_X1 U552 ( .A1(n518), .A2(n492), .ZN(n493) );
  XOR2_X1 U553 ( .A(G50GAT), .B(n493), .Z(G1331GAT) );
  NAND2_X1 U554 ( .A1(n564), .A2(n538), .ZN(n504) );
  OR2_X1 U555 ( .A1(n494), .A2(n504), .ZN(n499) );
  NOR2_X1 U556 ( .A1(n506), .A2(n499), .ZN(n495) );
  XOR2_X1 U557 ( .A(n495), .B(KEYINPUT42), .Z(n496) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(n496), .ZN(G1332GAT) );
  NOR2_X1 U559 ( .A1(n509), .A2(n499), .ZN(n497) );
  XOR2_X1 U560 ( .A(G64GAT), .B(n497), .Z(G1333GAT) );
  NOR2_X1 U561 ( .A1(n520), .A2(n499), .ZN(n498) );
  XOR2_X1 U562 ( .A(G71GAT), .B(n498), .Z(G1334GAT) );
  NOR2_X1 U563 ( .A1(n499), .A2(n518), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n501) );
  XNOR2_X1 U565 ( .A(G78GAT), .B(KEYINPUT103), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  OR2_X1 U568 ( .A1(n505), .A2(n504), .ZN(n512) );
  NOR2_X1 U569 ( .A1(n506), .A2(n512), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G85GAT), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n508), .B(n507), .ZN(G1336GAT) );
  NOR2_X1 U572 ( .A1(n509), .A2(n512), .ZN(n510) );
  XOR2_X1 U573 ( .A(G92GAT), .B(n510), .Z(G1337GAT) );
  NOR2_X1 U574 ( .A1(n520), .A2(n512), .ZN(n511) );
  XOR2_X1 U575 ( .A(G99GAT), .B(n511), .Z(G1338GAT) );
  NOR2_X1 U576 ( .A1(n518), .A2(n512), .ZN(n513) );
  XOR2_X1 U577 ( .A(KEYINPUT44), .B(n513), .Z(n514) );
  XNOR2_X1 U578 ( .A(G106GAT), .B(n514), .ZN(G1339GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(KEYINPUT109), .B(n517), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n518), .A2(n533), .ZN(n519) );
  NOR2_X1 U582 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U583 ( .A(KEYINPUT110), .B(n521), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n529), .A2(n535), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n524) );
  NAND2_X1 U587 ( .A1(n529), .A2(n538), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(G120GAT), .B(n525), .Z(G1341GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n527) );
  NAND2_X1 U591 ( .A1(n529), .A2(n543), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(G127GAT), .B(n528), .Z(G1342GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U595 ( .A1(n529), .A2(n547), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  XOR2_X1 U598 ( .A(G141GAT), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U599 ( .A1(n563), .A2(n533), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(n534), .Z(n548) );
  NAND2_X1 U601 ( .A1(n535), .A2(n548), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1344GAT) );
  XNOR2_X1 U603 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n542) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n540) );
  NAND2_X1 U605 ( .A1(n548), .A2(n538), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n545) );
  NAND2_X1 U609 ( .A1(n548), .A2(n543), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G155GAT), .B(n546), .ZN(G1346GAT) );
  XOR2_X1 U612 ( .A(G162GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n560), .A2(n564), .ZN(n552) );
  XNOR2_X1 U616 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n555) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(KEYINPUT56), .B(n556), .ZN(n559) );
  NOR2_X1 U623 ( .A1(n557), .A2(n560), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n571), .A2(n560), .ZN(n561) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n561), .Z(G1350GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n563), .ZN(n574) );
  NOR2_X1 U628 ( .A1(n564), .A2(n574), .ZN(n566) );
  XNOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  NOR2_X1 U632 ( .A1(n363), .A2(n574), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(G204GAT), .B(n570), .Z(G1353GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n574), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(n572), .Z(n573) );
  XNOR2_X1 U638 ( .A(G211GAT), .B(n573), .ZN(G1354GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

