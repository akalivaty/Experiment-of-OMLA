//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G57gat), .B(G64gat), .Z(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT97), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT97), .ZN(new_n212));
  XNOR2_X1  g011(.A(G71gat), .B(G78gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n205), .A2(new_n210), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT98), .ZN(new_n215));
  OR2_X1    g014(.A1(G57gat), .A2(G64gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G57gat), .A2(G64gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT95), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT95), .B1(new_n216), .B2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n206), .A2(KEYINPUT94), .ZN(new_n222));
  INV_X1    g021(.A(new_n206), .ZN(new_n223));
  INV_X1    g022(.A(G71gat), .ZN(new_n224));
  INV_X1    g023(.A(G78gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT94), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n222), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT96), .B1(new_n221), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT95), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n211), .B1(new_n232), .B2(new_n218), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT96), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(new_n234), .A3(new_n227), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n215), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT99), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(KEYINPUT99), .ZN(new_n241));
  INV_X1    g040(.A(G231gat), .ZN(new_n242));
  INV_X1    g041(.A(G233gat), .ZN(new_n243));
  NOR4_X1   g042(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n241), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n245), .A2(new_n239), .B1(G231gat), .B2(G233gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n204), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n245), .A2(G231gat), .A3(G233gat), .A4(new_n239), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n240), .A2(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n203), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n247), .B2(new_n250), .ZN(new_n255));
  XOR2_X1   g054(.A(G15gat), .B(G22gat), .Z(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT91), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT16), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(G1gat), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n257), .A2(G1gat), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(G8gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n236), .B2(new_n237), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n254), .A2(new_n255), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n250), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n251), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n268), .B2(new_n253), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n202), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n265), .B1(new_n254), .B2(new_n255), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n264), .A3(new_n253), .ZN(new_n272));
  INV_X1    g071(.A(new_n202), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G134gat), .B(G162gat), .Z(new_n276));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277));
  XOR2_X1   g076(.A(G43gat), .B(G50gat), .Z(new_n278));
  INV_X1    g077(.A(KEYINPUT15), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G43gat), .B(G50gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT15), .ZN(new_n282));
  NAND2_X1  g081(.A1(G29gat), .A2(G36gat), .ZN(new_n283));
  NOR3_X1   g082(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n280), .A2(new_n282), .A3(new_n283), .A4(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n286), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n284), .B1(new_n289), .B2(KEYINPUT89), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT89), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n290), .A2(new_n292), .B1(G29gat), .B2(G36gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n293), .B2(new_n282), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT90), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n294), .A2(new_n299), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n302));
  NAND2_X1  g101(.A1(G85gat), .A2(G92gat), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(G85gat), .A2(G92gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n302), .B2(new_n303), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G99gat), .B(G106gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT101), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n309), .A2(G99gat), .A3(G106gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(G99gat), .B2(G106gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT8), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n307), .A2(KEYINPUT102), .A3(new_n308), .A4(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n304), .A2(new_n306), .A3(new_n312), .A4(new_n308), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT102), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n304), .A2(new_n312), .A3(new_n306), .ZN(new_n317));
  INV_X1    g116(.A(new_n308), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n300), .A2(new_n301), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n296), .A2(new_n297), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT41), .ZN(new_n324));
  INV_X1    g123(.A(G232gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n243), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OAI22_X1  g126(.A1(new_n323), .A2(new_n320), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n277), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n324), .ZN(new_n330));
  INV_X1    g129(.A(new_n328), .ZN(new_n331));
  INV_X1    g130(.A(new_n277), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n321), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n329), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n330), .B1(new_n329), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n276), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  INV_X1    g137(.A(new_n276), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n334), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n298), .A2(new_n262), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n262), .B1(new_n296), .B2(new_n297), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G229gat), .A2(G233gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT13), .Z(new_n348));
  AOI21_X1  g147(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n323), .A2(new_n263), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n342), .B(new_n348), .C1(new_n350), .C2(new_n344), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n323), .A2(KEYINPUT17), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n263), .A2(new_n301), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n343), .B(new_n347), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT18), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n300), .A2(new_n263), .A3(new_n301), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n359), .A2(KEYINPUT18), .A3(new_n347), .A4(new_n343), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G113gat), .B(G141gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT11), .ZN(new_n363));
  INV_X1    g162(.A(G169gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G197gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT12), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT93), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n358), .B(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n360), .B(new_n368), .C1(new_n349), .C2(new_n352), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n361), .A2(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n236), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n314), .A3(new_n319), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT103), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n320), .A2(new_n236), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n320), .B2(new_n236), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n377), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n320), .A2(new_n236), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G230gat), .A2(G233gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n388));
  INV_X1    g187(.A(new_n386), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G120gat), .B(G148gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G176gat), .B(G204gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n275), .A2(new_n341), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n402));
  NOR2_X1   g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G169gat), .A2(G176gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT26), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(KEYINPUT26), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT27), .B(G183gat), .ZN(new_n412));
  INV_X1    g211(.A(G190gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(new_n413), .C1(KEYINPUT67), .C2(KEYINPUT28), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT66), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT25), .ZN(new_n421));
  NAND3_X1  g220(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n424), .A2(new_n425), .B1(new_n410), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n403), .A2(KEYINPUT23), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT23), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(G169gat), .B2(G176gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n430), .B2(new_n403), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n420), .B(new_n421), .C1(new_n427), .C2(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n429), .A2(G169gat), .A3(G176gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n405), .A2(KEYINPUT23), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n404), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(new_n410), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n422), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(KEYINPUT25), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n425), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n436), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n435), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n420), .B1(new_n442), .B2(new_n421), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n419), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT68), .B(G120gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G113gat), .ZN(new_n446));
  INV_X1    g245(.A(G120gat), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT69), .B1(new_n447), .B2(G113gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n449));
  INV_X1    g248(.A(G113gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(G120gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G127gat), .B(G134gat), .Z(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT1), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT1), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n447), .A2(G113gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n450), .A2(G120gat), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n453), .A2(new_n455), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT64), .Z(new_n463));
  INV_X1    g262(.A(new_n460), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n419), .B(new_n464), .C1(new_n439), .C2(new_n443), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(KEYINPUT32), .ZN(new_n469));
  XOR2_X1   g268(.A(G15gat), .B(G43gat), .Z(new_n470));
  XNOR2_X1  g269(.A(G71gat), .B(G99gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n466), .B(KEYINPUT32), .C1(new_n467), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n463), .B1(new_n461), .B2(new_n465), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n479));
  NOR3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n479), .ZN(new_n481));
  INV_X1    g280(.A(new_n463), .ZN(new_n482));
  INV_X1    g281(.A(new_n465), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n421), .B1(new_n427), .B2(new_n431), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT66), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n432), .A3(new_n438), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n464), .B1(new_n486), .B2(new_n419), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n482), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n488), .B2(KEYINPUT70), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n476), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n479), .B1(new_n477), .B2(new_n478), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(KEYINPUT70), .A3(new_n481), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n475), .B2(new_n473), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT86), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G78gat), .B(G106gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n497), .B(KEYINPUT79), .Z(new_n498));
  AND2_X1   g297(.A1(G155gat), .A2(G162gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(G155gat), .A2(G162gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT77), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G155gat), .ZN(new_n502));
  INV_X1    g301(.A(G162gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT77), .ZN(new_n505));
  NAND2_X1  g304(.A1(G155gat), .A2(G162gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(KEYINPUT2), .ZN(new_n509));
  INV_X1    g308(.A(G148gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G141gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G141gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G148gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n508), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT75), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT74), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n506), .A2(new_n520), .A3(KEYINPUT2), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G141gat), .B(G148gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n506), .B2(KEYINPUT2), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT73), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G155gat), .B2(G162gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n506), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(KEYINPUT73), .B2(new_n506), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n519), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n511), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n506), .B2(new_n527), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(KEYINPUT75), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n518), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G197gat), .B(G204gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  XNOR2_X1  g338(.A(G211gat), .B(G218gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G211gat), .ZN(new_n543));
  INV_X1    g342(.A(G218gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n540), .B(new_n538), .C1(KEYINPUT22), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT3), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT82), .B1(new_n537), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT3), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n508), .A2(new_n509), .A3(new_n517), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n533), .A2(KEYINPUT75), .A3(new_n535), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT75), .B1(new_n533), .B2(new_n535), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT82), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n542), .A2(KEYINPUT72), .A3(new_n546), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT72), .B1(new_n542), .B2(new_n546), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n552), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n566), .B2(KEYINPUT29), .ZN(new_n567));
  NAND2_X1  g366(.A1(G228gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n560), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(KEYINPUT80), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT81), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n546), .B1(new_n542), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT81), .B1(new_n539), .B2(new_n541), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n548), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n537), .B1(new_n552), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n563), .B1(new_n565), .B2(new_n548), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G22gat), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n570), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n498), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n570), .A2(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G22gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n585));
  INV_X1    g384(.A(new_n498), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G50gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n582), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n580), .A2(new_n581), .A3(new_n498), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n586), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n476), .A2(new_n490), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT86), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n494), .A2(new_n475), .A3(new_n473), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n496), .A2(new_n590), .A3(new_n594), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G1gat), .B(G29gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT0), .ZN(new_n601));
  XNOR2_X1  g400(.A(G57gat), .B(G85gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n557), .A2(KEYINPUT3), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n464), .A3(new_n565), .ZN(new_n605));
  NAND2_X1  g404(.A1(G225gat), .A2(G233gat), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n460), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT4), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n537), .A2(KEYINPUT4), .A3(new_n460), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n605), .A2(new_n606), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT5), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n606), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n537), .A2(new_n460), .ZN(new_n616));
  INV_X1    g415(.A(new_n607), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n612), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n603), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n464), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n530), .A2(new_n536), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n552), .B1(new_n622), .B2(new_n554), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n609), .B(new_n610), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n618), .B1(new_n624), .B2(new_n615), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT5), .ZN(new_n626));
  INV_X1    g425(.A(new_n603), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n613), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT6), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n626), .A2(KEYINPUT6), .A3(new_n627), .A4(new_n613), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G8gat), .B(G36gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G64gat), .B(G92gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G226gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n243), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n419), .B(new_n637), .C1(new_n439), .C2(new_n443), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n548), .B1(new_n636), .B2(new_n243), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n486), .B2(new_n419), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n564), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n432), .A2(new_n438), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n643), .A2(new_n485), .B1(new_n418), .B2(new_n411), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n638), .B(new_n563), .C1(new_n644), .C2(new_n640), .ZN(new_n645));
  AOI211_X1 g444(.A(KEYINPUT30), .B(new_n635), .C1(new_n642), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT30), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n645), .ZN(new_n648));
  INV_X1    g447(.A(new_n635), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n645), .A3(new_n635), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n632), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n402), .B1(new_n599), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n654), .B(new_n652), .C1(new_n630), .C2(new_n631), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n582), .A2(new_n587), .A3(new_n589), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n589), .B1(new_n582), .B2(new_n587), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n660), .A2(new_n661), .A3(KEYINPUT88), .A4(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n491), .A2(new_n495), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n594), .A3(new_n590), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n632), .A2(new_n653), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT35), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n657), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n666), .B(KEYINPUT36), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n594), .A2(new_n590), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT37), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT84), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT37), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n648), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n649), .A2(KEYINPUT38), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n674), .B2(KEYINPUT84), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT85), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n635), .B1(new_n642), .B2(new_n645), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n674), .A3(new_n635), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(KEYINPUT38), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n679), .A2(KEYINPUT85), .A3(new_n681), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n632), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n624), .A2(new_n615), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT39), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n616), .A2(new_n617), .A3(new_n615), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(new_n690), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n691), .B(new_n603), .C1(new_n689), .C2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(KEYINPUT83), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n693), .A2(new_n689), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(KEYINPUT83), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n697), .A2(new_n603), .A3(new_n691), .A4(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n696), .A2(new_n628), .A3(new_n652), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n664), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n671), .B(new_n673), .C1(new_n688), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n670), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n401), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n632), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT105), .B(G1gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1324gat));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n653), .ZN(new_n708));
  INV_X1    g507(.A(G8gat), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  MUX2_X1   g511(.A(KEYINPUT42), .B(new_n710), .S(new_n712), .Z(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n704), .B2(new_n671), .ZN(new_n714));
  INV_X1    g513(.A(new_n660), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(G15gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n704), .B2(new_n716), .ZN(G1326gat));
  NOR2_X1   g516(.A1(new_n704), .A2(new_n664), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n341), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n337), .A2(new_n340), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n670), .B2(new_n702), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n275), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n400), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n721), .B1(new_n732), .B2(new_n632), .ZN(new_n733));
  INV_X1    g532(.A(new_n632), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(G29gat), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n730), .A2(new_n726), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(G29gat), .A3(new_n632), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT45), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(G1328gat));
  OAI21_X1  g539(.A(G36gat), .B1(new_n732), .B2(new_n653), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n737), .A2(G36gat), .A3(new_n653), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1329gat));
  INV_X1    g543(.A(new_n671), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n731), .A2(G43gat), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n737), .A2(new_n715), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(G43gat), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g548(.A1(new_n731), .A2(G50gat), .A3(new_n672), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n737), .A2(new_n664), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(G50gat), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1331gat));
  NAND4_X1  g553(.A1(new_n270), .A2(new_n725), .A3(new_n274), .A4(new_n374), .ZN(new_n755));
  AOI211_X1 g554(.A(new_n399), .B(new_n755), .C1(new_n702), .C2(new_n670), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n734), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g557(.A(new_n653), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT108), .Z(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n761), .B(new_n762), .Z(G1333gat));
  XOR2_X1   g562(.A(new_n660), .B(KEYINPUT109), .Z(new_n764));
  AOI21_X1  g563(.A(G71gat), .B1(new_n756), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n671), .A2(new_n224), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n756), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g567(.A1(new_n756), .A2(new_n672), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  INV_X1    g569(.A(G85gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n275), .A2(new_n374), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n399), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n724), .A2(new_n727), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT110), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n724), .A2(new_n776), .A3(new_n727), .A4(new_n773), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n734), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n771), .B1(new_n778), .B2(KEYINPUT111), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(KEYINPUT111), .B2(new_n778), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n722), .B2(new_n772), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n726), .A2(KEYINPUT51), .A3(new_n275), .A4(new_n374), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n734), .A2(new_n771), .A3(new_n398), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(G1336gat));
  NAND3_X1  g586(.A1(new_n775), .A2(new_n652), .A3(new_n777), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(KEYINPUT112), .A3(new_n783), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n399), .A2(G92gat), .A3(new_n653), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n781), .C1(new_n722), .C2(new_n772), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(new_n792), .A3(new_n794), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n789), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT114), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT52), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(new_n784), .B2(new_n792), .ZN(new_n803));
  OAI21_X1  g602(.A(G92gat), .B1(new_n774), .B2(new_n653), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(new_n802), .A3(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n775), .A2(new_n745), .A3(new_n777), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n715), .A2(G99gat), .A3(new_n399), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n785), .B2(new_n809), .ZN(G1338gat));
  NAND3_X1  g609(.A1(new_n775), .A2(new_n672), .A3(new_n777), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n790), .A2(new_n794), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n399), .A2(new_n664), .A3(G106gat), .ZN(new_n813));
  AOI22_X1  g612(.A1(G106gat), .A2(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n784), .B2(new_n813), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  OAI21_X1  g616(.A(G106gat), .B1(new_n774), .B2(new_n664), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n816), .B2(new_n818), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n814), .A2(new_n815), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NOR2_X1   g620(.A1(new_n632), .A2(new_n652), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n382), .A2(new_n384), .A3(new_n389), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n387), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n389), .B1(new_n382), .B2(new_n384), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n396), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n374), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n829), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n826), .A2(new_n829), .A3(new_n834), .A4(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT117), .B1(new_n836), .B2(new_n397), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838));
  INV_X1    g637(.A(new_n397), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n838), .B(new_n839), .C1(new_n833), .C2(new_n835), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n831), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n359), .A2(new_n343), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(G229gat), .A3(G233gat), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n346), .A2(new_n348), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n367), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n371), .B2(new_n373), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n398), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT118), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n341), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n837), .A2(new_n840), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n830), .A2(new_n824), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n341), .A2(new_n851), .A3(new_n846), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n275), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n755), .A2(new_n398), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n667), .B(new_n823), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n375), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n599), .B(new_n823), .C1(new_n854), .C2(new_n855), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n374), .A2(new_n450), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n445), .A3(new_n398), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n854), .A2(new_n855), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n822), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n599), .A3(new_n399), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n864), .B2(new_n447), .ZN(G1341gat));
  NAND2_X1  g664(.A1(new_n858), .A2(new_n729), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n275), .A2(G127gat), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n866), .A2(G127gat), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT119), .ZN(G1342gat));
  NOR4_X1   g668(.A1(new_n863), .A2(G134gat), .A3(new_n667), .A4(new_n725), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT56), .ZN(new_n871));
  INV_X1    g670(.A(G134gat), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n863), .A2(new_n599), .A3(new_n725), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n745), .A2(new_n823), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n862), .B2(new_n672), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n672), .A2(KEYINPUT57), .ZN(new_n877));
  INV_X1    g676(.A(new_n853), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n375), .A2(new_n851), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n836), .A2(new_n397), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n847), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n725), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n275), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n877), .B1(new_n884), .B2(new_n855), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n375), .B(new_n875), .C1(new_n876), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n745), .A2(new_n664), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n374), .A2(G141gat), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n862), .A2(new_n822), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n890), .B(KEYINPUT120), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1344gat));
  NOR4_X1   g695(.A1(new_n399), .A2(G148gat), .A3(new_n632), .A4(new_n652), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n862), .A2(new_n888), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n875), .B1(new_n876), .B2(new_n885), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n399), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(KEYINPUT59), .A3(new_n510), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n862), .A2(new_n672), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n664), .A2(KEYINPUT57), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n729), .B1(new_n878), .B2(new_n882), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n755), .A2(new_n907), .A3(new_n398), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n755), .B2(new_n398), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n904), .A2(new_n398), .A3(new_n875), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n902), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n898), .B1(new_n901), .B2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n899), .B2(new_n275), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n863), .A2(new_n664), .A3(new_n745), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n502), .A3(new_n729), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1346gat));
  OAI211_X1 g717(.A(new_n341), .B(new_n875), .C1(new_n876), .C2(new_n885), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G162gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n503), .A3(new_n341), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n734), .A2(new_n653), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n862), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n667), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n375), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n764), .A2(new_n664), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(new_n364), .A3(new_n374), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n931), .A2(new_n934), .ZN(G1348gat));
  INV_X1    g734(.A(G176gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n936), .A3(new_n398), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n933), .B2(new_n399), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n933), .B2(new_n275), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n928), .A2(new_n412), .A3(new_n929), .A4(new_n729), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n341), .A3(new_n932), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n948), .A3(G190gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n947), .A2(new_n951), .A3(new_n948), .A4(G190gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n947), .A2(G190gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n930), .A2(new_n413), .A3(new_n341), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1351gat));
  NAND3_X1  g756(.A1(new_n928), .A2(KEYINPUT125), .A3(new_n888), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n862), .A2(new_n888), .A3(new_n927), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n958), .A2(new_n366), .A3(new_n375), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n671), .A2(new_n927), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n664), .B1(new_n854), .B2(new_n855), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT57), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n911), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n374), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n962), .A2(new_n971), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n959), .A2(G204gat), .A3(new_n399), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n904), .A2(new_n398), .A3(new_n911), .ZN(new_n976));
  OAI21_X1  g775(.A(G204gat), .B1(new_n976), .B2(new_n963), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1353gat));
  OAI211_X1 g777(.A(KEYINPUT63), .B(G211gat), .C1(new_n967), .C2(new_n275), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n904), .A2(new_n729), .A3(new_n911), .A4(new_n964), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(G211gat), .B1(new_n967), .B2(new_n275), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT63), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n980), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n958), .A2(new_n543), .A3(new_n729), .A4(new_n961), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n967), .B2(new_n725), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n958), .A2(new_n961), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n341), .A2(new_n544), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G1355gat));
endmodule


