//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n594, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND2_X1  g026(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT70), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT71), .A3(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT72), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n483), .A3(G101), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n479), .A2(G2105), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n469), .B1(new_n465), .B2(new_n467), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n473), .A2(G136), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n469), .A2(G138), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n476), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT3), .B1(new_n466), .B2(G2104), .ZN(new_n501));
  OAI211_X1 g076(.A(KEYINPUT73), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n465), .B2(new_n467), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT73), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n469), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n491), .B2(G126), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(KEYINPUT74), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT74), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT75), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n526), .B1(new_n523), .B2(KEYINPUT75), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n517), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT6), .B1(new_n514), .B2(new_n515), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n520), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n522), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n531), .B2(new_n533), .ZN(new_n538));
  AOI22_X1  g113(.A1(G50), .A2(new_n534), .B1(new_n538), .B2(G88), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n528), .A2(new_n529), .ZN(new_n541));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n528), .A2(new_n529), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n543), .A2(new_n530), .A3(new_n544), .A4(new_n539), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G166));
  NAND2_X1  g121(.A1(new_n534), .A2(G51), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n521), .A2(new_n522), .ZN(new_n551));
  AND2_X1   g126(.A1(G63), .A2(G651), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n549), .A2(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n538), .A2(G89), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(G286));
  INV_X1    g131(.A(G286), .ZN(G168));
  AOI22_X1  g132(.A1(new_n551), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n516), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT78), .ZN(new_n560));
  AOI22_X1  g135(.A1(G52), .A2(new_n534), .B1(new_n538), .B2(G90), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G171));
  AOI22_X1  g138(.A1(new_n551), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n516), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(G43), .B2(new_n534), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n538), .A2(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT80), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n537), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n538), .A2(G91), .B1(new_n579), .B2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n582));
  INV_X1    g157(.A(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n581), .B1(new_n584), .B2(new_n513), .ZN(new_n585));
  OAI211_X1 g160(.A(G53), .B(G543), .C1(new_n585), .C2(new_n532), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n580), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(G299));
  NAND2_X1  g166(.A1(new_n562), .A2(KEYINPUT82), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n562), .A2(KEYINPUT82), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(G301));
  INV_X1    g170(.A(G166), .ZN(G303));
  NAND2_X1  g171(.A1(new_n534), .A2(G49), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n538), .A2(G87), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n551), .B2(G74), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n521), .B2(new_n522), .ZN(new_n602));
  AND2_X1   g177(.A1(G73), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n517), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g179(.A(G48), .B(G543), .C1(new_n585), .C2(new_n532), .ZN(new_n605));
  OAI211_X1 g180(.A(G86), .B(new_n551), .C1(new_n585), .C2(new_n532), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(new_n534), .A2(G47), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n538), .A2(G85), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT84), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n551), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n516), .B1(new_n612), .B2(KEYINPUT83), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT83), .B2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(new_n538), .A2(G92), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT10), .Z(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n537), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n534), .A2(G54), .B1(new_n620), .B2(G651), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n622), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g198(.A(new_n622), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n589), .B(KEYINPUT81), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(new_n622), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n569), .ZN(G323));
  XOR2_X1   g209(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n635));
  XNOR2_X1  g210(.A(G323), .B(new_n635), .ZN(G282));
  NAND2_X1  g211(.A1(new_n476), .A2(new_n480), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT13), .B(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n473), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n491), .A2(G123), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(G2096), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT88), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2451), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n654), .B(new_n660), .Z(new_n661));
  XOR2_X1   g236(.A(KEYINPUT87), .B(KEYINPUT16), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2454), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(G14), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n661), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  INV_X1    g247(.A(new_n669), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n673), .B2(new_n667), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n667), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n674), .B1(new_n677), .B2(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n673), .A3(new_n670), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n685), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  NAND2_X1  g279(.A1(new_n629), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G4), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G32), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n713), .A2(new_n714), .B1(G105), .B2(new_n480), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n473), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n491), .A2(G129), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n710), .B1(new_n719), .B2(new_n709), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT27), .B(G1996), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT97), .B(G2067), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n709), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n491), .A2(G128), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n473), .A2(G140), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n469), .A2(G116), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n722), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n723), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n720), .A2(new_n721), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G28), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n709), .B1(new_n736), .B2(G28), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n735), .B1(new_n737), .B2(new_n738), .C1(new_n646), .C2(new_n709), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G19), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n569), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G1341), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n734), .B(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n706), .A2(new_n707), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n708), .A2(new_n733), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n709), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n709), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT29), .Z(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G2090), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n709), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  NOR2_X1   g328(.A1(G27), .A2(G29), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n750), .A2(G2090), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n746), .A2(new_n751), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G5), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G171), .B2(new_n760), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT24), .B(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(new_n709), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT99), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n486), .B2(new_n709), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n762), .A2(G1961), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(new_n743), .B2(new_n742), .C1(G1961), .C2(new_n762), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n760), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n760), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT100), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G1966), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n709), .A2(G33), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n476), .A2(G127), .ZN(new_n775));
  INV_X1    g350(.A(G115), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n464), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n469), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(new_n473), .B2(G139), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n774), .B1(new_n787), .B2(new_n709), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G2072), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G2072), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n789), .B(new_n790), .C1(new_n763), .C2(new_n767), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n769), .A2(new_n773), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n772), .A2(G1966), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT101), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n760), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n626), .B2(new_n760), .ZN(new_n797));
  INV_X1    g372(.A(G1956), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n759), .A2(new_n792), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n760), .A2(G23), .ZN(new_n801));
  INV_X1    g376(.A(G288), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n760), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT33), .ZN(new_n804));
  INV_X1    g379(.A(G1976), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n760), .A2(G6), .ZN(new_n807));
  INV_X1    g382(.A(G305), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n760), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT32), .B(G1981), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT94), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT95), .Z(new_n813));
  NOR2_X1   g388(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n815));
  NAND2_X1  g390(.A1(G166), .A2(G16), .ZN(new_n816));
  NOR2_X1   g391(.A1(G16), .A2(G22), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g394(.A(KEYINPUT96), .B(new_n817), .C1(G166), .C2(G16), .ZN(new_n820));
  INV_X1    g395(.A(G1971), .ZN(new_n821));
  OR3_X1    g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n819), .B2(new_n820), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n814), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n760), .A2(G24), .ZN(new_n827));
  INV_X1    g402(.A(G290), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n760), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1986), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n709), .A2(G25), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT92), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n491), .A2(G119), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n473), .A2(G131), .ZN(new_n834));
  OR2_X1    g409(.A1(G95), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT93), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n832), .B1(new_n839), .B2(G29), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G1991), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n830), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n825), .A2(new_n826), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n825), .A2(new_n846), .A3(new_n826), .A4(new_n843), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n800), .B1(new_n845), .B2(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n847), .ZN(new_n849));
  INV_X1    g424(.A(new_n800), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(G150));
  NAND2_X1  g426(.A1(new_n629), .A2(G559), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n538), .A2(G93), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n534), .A2(G55), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n551), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n854), .B(new_n855), .C1(new_n516), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n568), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(KEYINPUT39), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT102), .B(G860), .Z(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(G145));
  XOR2_X1   g442(.A(new_n511), .B(KEYINPUT103), .Z(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n473), .A2(G142), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n491), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n469), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n837), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n639), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n834), .A2(new_n833), .A3(new_n836), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n639), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n787), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n719), .B(new_n730), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n786), .A3(new_n880), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n869), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n868), .A3(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n494), .B(new_n646), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G160), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  INV_X1    g471(.A(new_n894), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n888), .A2(new_n890), .A3(new_n891), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n896), .A4(new_n898), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT40), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(G395));
  INV_X1    g480(.A(G868), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n857), .A2(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n858), .B(KEYINPUT106), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n632), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n626), .A2(KEYINPUT107), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n629), .ZN(new_n913));
  NAND3_X1  g488(.A1(G299), .A2(new_n910), .A3(new_n622), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n914), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(G303), .A2(G305), .ZN(new_n921));
  NAND2_X1  g496(.A1(G166), .A2(new_n808), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n802), .B1(new_n611), .B2(new_n614), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n611), .A2(new_n802), .A3(new_n614), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n923), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT108), .B1(new_n929), .B2(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n924), .A3(new_n927), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n921), .A4(new_n922), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n933), .B2(new_n936), .ZN(new_n938));
  OAI221_X1 g513(.A(new_n916), .B1(new_n909), .B2(new_n920), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n916), .B1(new_n909), .B2(new_n920), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n907), .B1(new_n943), .B2(new_n906), .ZN(G295));
  OAI21_X1  g519(.A(new_n907), .B1(new_n943), .B2(new_n906), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n946), .B2(KEYINPUT110), .ZN(new_n947));
  INV_X1    g522(.A(new_n858), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT82), .ZN(new_n949));
  NAND2_X1  g524(.A1(G171), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G286), .B1(new_n950), .B2(new_n592), .ZN(new_n951));
  NOR2_X1   g526(.A1(G171), .A2(G168), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n952), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n858), .B(new_n954), .C1(G301), .C2(G286), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n918), .A2(new_n919), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n955), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n914), .A3(new_n913), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n933), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n958), .A3(new_n932), .A4(new_n928), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(new_n946), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n946), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n947), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n933), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n896), .A3(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n946), .A3(new_n961), .ZN(new_n968));
  INV_X1    g543(.A(new_n947), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n970), .ZN(G397));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(G1384), .ZN(new_n972));
  INV_X1    g547(.A(new_n499), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n496), .B1(new_n504), .B2(KEYINPUT73), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT73), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n510), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT45), .B(new_n972), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n475), .A2(new_n485), .A3(G40), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n506), .B2(new_n510), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n980), .B(new_n981), .C1(new_n982), .C2(KEYINPUT45), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n475), .A2(new_n485), .A3(G40), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n978), .B2(new_n979), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(KEYINPUT113), .A3(new_n980), .ZN(new_n991));
  AOI21_X1  g566(.A(G2078), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(KEYINPUT53), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n982), .A2(KEYINPUT45), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n753), .A2(KEYINPUT53), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n990), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n986), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(new_n987), .C1(new_n978), .C2(new_n979), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1961), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT122), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n981), .B1(new_n982), .B2(new_n999), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1000), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n996), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(G301), .B1(new_n993), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n605), .A2(new_n604), .A3(new_n606), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT116), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n981), .A2(new_n982), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n597), .A2(new_n598), .A3(G1976), .A4(new_n599), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT115), .Z(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n805), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n1016), .A4(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1022), .B(KEYINPUT115), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1021), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n985), .A2(new_n991), .A3(new_n821), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT114), .B(G2090), .Z(new_n1031));
  NAND3_X1  g606(.A1(new_n998), .A2(new_n1000), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n542), .A2(G8), .A3(new_n545), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n542), .A2(new_n545), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1028), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n982), .A2(KEYINPUT117), .A3(new_n999), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1000), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n998), .A3(new_n1031), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1030), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1038), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1010), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1966), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n981), .B1(new_n982), .B2(KEYINPUT45), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n988), .A2(new_n989), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n998), .A2(new_n763), .A3(new_n1000), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G168), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(G168), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT51), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1060), .A3(G8), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT126), .B1(new_n1049), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1038), .A3(G8), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1028), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1038), .B1(G8), .B2(new_n1045), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1010), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(new_n1059), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1063), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1021), .A2(new_n805), .A3(new_n802), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1013), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1018), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1065), .B2(new_n1028), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1039), .A2(new_n1048), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1082), .A2(new_n1029), .A3(G286), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1039), .A2(new_n1086), .A3(KEYINPUT63), .A4(new_n1083), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1079), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1956), .B1(new_n1043), .B2(new_n998), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n988), .A2(new_n989), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT56), .B(G2072), .Z(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(new_n981), .A3(new_n980), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n580), .B(new_n1095), .C1(new_n587), .C2(new_n588), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n586), .B(KEYINPUT9), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1098), .B2(new_n580), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1089), .A2(new_n1094), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT117), .B1(new_n982), .B2(new_n999), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1000), .A2(new_n1041), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n998), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n798), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1100), .B1(new_n1106), .B2(new_n1093), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1348), .B1(new_n998), .B2(new_n1000), .ZN(new_n1108));
  INV_X1    g683(.A(G2067), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n981), .A2(new_n982), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n629), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1102), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1093), .A2(new_n1100), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1106), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1101), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n988), .B2(new_n986), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n983), .B2(G1996), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n569), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(new_n569), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1119), .A2(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1117), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT120), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n707), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT60), .B1(new_n1133), .B2(new_n1110), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1134), .A2(KEYINPUT121), .A3(new_n622), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1138), .B2(new_n629), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1132), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT121), .B1(new_n1134), .B2(new_n622), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1136), .A3(new_n629), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1142), .A4(new_n1131), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1130), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT120), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1116), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1008), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1007), .B1(new_n1006), .B2(new_n996), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(new_n992), .B2(KEYINPUT53), .ZN(new_n1150));
  INV_X1    g725(.A(G301), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n511), .A2(new_n972), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n989), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT53), .B1(new_n1156), .B2(G2078), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n1156), .B2(G2078), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n980), .A2(new_n981), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1001), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n993), .A2(new_n1153), .A3(G301), .A4(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1160), .B(G301), .C1(new_n992), .C2(KEYINPUT53), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT124), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1152), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n993), .A2(new_n1160), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1167), .B2(G171), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT125), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n993), .A2(new_n1009), .A3(new_n1170), .A4(G301), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1081), .A2(new_n1073), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1166), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1075), .B(new_n1088), .C1(new_n1147), .C2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1155), .A2(new_n986), .ZN(new_n1176));
  INV_X1    g751(.A(G1986), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n828), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT112), .Z(new_n1179));
  XNOR2_X1  g754(.A(new_n730), .B(new_n1109), .ZN(new_n1180));
  INV_X1    g755(.A(G1996), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n718), .B(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n878), .B(new_n841), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1183), .B(new_n1184), .C1(new_n828), .C2(new_n1177), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1176), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1175), .A2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1179), .A2(new_n1176), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1188), .A2(KEYINPUT48), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1179), .A2(KEYINPUT48), .A3(new_n1176), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1176), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1180), .A2(new_n719), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1195), .A2(new_n1196), .B1(new_n1176), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT47), .Z(new_n1199));
  NAND2_X1  g774(.A1(new_n838), .A2(new_n841), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT127), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1183), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1200), .A2(KEYINPUT127), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1202), .A2(new_n1203), .B1(G2067), .B2(new_n730), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1176), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1193), .A2(new_n1199), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1187), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g782(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n703), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n901), .B2(new_n902), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n968), .ZN(new_n1212));
  AND2_X1   g786(.A1(new_n1211), .A2(new_n1212), .ZN(G308));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(G225));
endmodule


