//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1109, new_n1110,
    new_n1111, new_n1113, new_n1114, new_n1115, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179;
  NOR2_X1   g000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g001(.A(G50), .ZN(new_n202));
  NAND2_X1  g002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g005(.A(G1), .ZN(new_n206));
  INV_X1    g006(.A(G20), .ZN(new_n207));
  NOR2_X1   g007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  OAI21_X1  g015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g017(.A(G58), .ZN(new_n218));
  INV_X1    g018(.A(G232), .ZN(new_n219));
  INV_X1    g019(.A(G107), .ZN(new_n220));
  INV_X1    g020(.A(G264), .ZN(new_n221));
  OAI221_X1 g021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g029(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  XNOR2_X1  g033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g036(.A(new_n236), .B(new_n219), .ZN(new_n237));
  XOR2_X1   g037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g047(.A(G13), .ZN(new_n248));
  NOR3_X1   g048(.A1(new_n248), .A2(new_n207), .A3(G1), .ZN(new_n249));
  NAND3_X1  g049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n213), .ZN(new_n251));
  NOR2_X1   g051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g052(.A1(new_n206), .A2(G20), .ZN(new_n253));
  NAND3_X1  g053(.A1(new_n252), .A2(G50), .A3(new_n253), .ZN(new_n254));
  INV_X1    g054(.A(new_n249), .ZN(new_n255));
  OAI21_X1  g055(.A(new_n254), .B1(G50), .B2(new_n255), .ZN(new_n256));
  INV_X1    g056(.A(G33), .ZN(new_n257));
  NAND2_X1  g057(.A1(new_n207), .A2(new_n257), .ZN(new_n258));
  INV_X1    g058(.A(new_n258), .ZN(new_n259));
  AOI22_X1  g059(.A1(G150), .A2(new_n259), .B1(new_n203), .B2(G20), .ZN(new_n260));
  NAND2_X1  g060(.A1(new_n207), .A2(G33), .ZN(new_n261));
  XNOR2_X1  g061(.A(new_n261), .B(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  OAI21_X1  g063(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g064(.A(new_n256), .B1(new_n251), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g065(.A(new_n265), .B(KEYINPUT9), .Z(new_n266));
  INV_X1    g066(.A(G41), .ZN(new_n267));
  NOR2_X1   g067(.A1(new_n257), .A2(new_n267), .ZN(new_n268));
  MUX2_X1   g068(.A(G222), .B(G223), .S(G1698), .Z(new_n269));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g071(.A(G77), .ZN(new_n272));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n270), .ZN(new_n273));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n274));
  AOI211_X1 g074(.A(new_n213), .B(new_n268), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  OAI21_X1  g075(.A(new_n275), .B1(new_n274), .B2(new_n273), .ZN(new_n276));
  AOI21_X1  g076(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g077(.A(G274), .ZN(new_n278));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g079(.A(KEYINPUT66), .B(G41), .ZN(new_n280));
  INV_X1    g080(.A(G45), .ZN(new_n281));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g082(.A1(new_n279), .A2(new_n206), .A3(new_n282), .ZN(new_n283));
  INV_X1    g083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g084(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n285));
  OAI21_X1  g085(.A(new_n285), .B1(new_n268), .B2(new_n213), .ZN(new_n286));
  XNOR2_X1  g086(.A(new_n286), .B(KEYINPUT67), .ZN(new_n287));
  AOI21_X1  g087(.A(new_n284), .B1(new_n287), .B2(G226), .ZN(new_n288));
  NAND2_X1  g088(.A1(new_n276), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  INV_X1    g090(.A(G190), .ZN(new_n291));
  OAI211_X1 g091(.A(new_n266), .B(new_n290), .C1(new_n291), .C2(new_n289), .ZN(new_n292));
  XNOR2_X1  g092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g093(.A(G169), .ZN(new_n294));
  AOI21_X1  g094(.A(new_n265), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g095(.A(new_n295), .B1(G179), .B2(new_n289), .ZN(new_n296));
  AND2_X1   g096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g097(.A1(new_n287), .A2(G244), .ZN(new_n298));
  INV_X1    g098(.A(G1698), .ZN(new_n299));
  NAND2_X1  g099(.A1(new_n270), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g100(.A(KEYINPUT70), .B(G107), .ZN(new_n301));
  INV_X1    g101(.A(new_n301), .ZN(new_n302));
  OAI22_X1  g102(.A1(new_n300), .A2(new_n219), .B1(new_n302), .B2(new_n270), .ZN(new_n303));
  NAND2_X1  g103(.A1(new_n270), .A2(G1698), .ZN(new_n304));
  INV_X1    g104(.A(G238), .ZN(new_n305));
  NOR2_X1   g105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g106(.A(new_n277), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g107(.A1(new_n298), .A2(new_n283), .A3(new_n307), .ZN(new_n308));
  INV_X1    g108(.A(new_n308), .ZN(new_n309));
  INV_X1    g109(.A(G179), .ZN(new_n310));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g111(.A(new_n251), .ZN(new_n312));
  INV_X1    g112(.A(new_n263), .ZN(new_n313));
  AOI22_X1  g113(.A1(new_n313), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n314));
  XNOR2_X1  g114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  OR2_X1    g115(.A1(new_n262), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g116(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g117(.A1(new_n252), .A2(G77), .A3(new_n253), .ZN(new_n318));
  OAI21_X1  g118(.A(new_n318), .B1(G77), .B2(new_n255), .ZN(new_n319));
  NOR2_X1   g119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g121(.A1(new_n308), .A2(new_n294), .ZN(new_n322));
  NAND3_X1  g122(.A1(new_n311), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g123(.A(G200), .ZN(new_n324));
  OAI21_X1  g124(.A(new_n320), .B1(new_n309), .B2(new_n324), .ZN(new_n325));
  AOI22_X1  g125(.A1(new_n325), .A2(KEYINPUT71), .B1(G190), .B2(new_n309), .ZN(new_n326));
  OAI21_X1  g126(.A(new_n326), .B1(KEYINPUT71), .B2(new_n325), .ZN(new_n327));
  NAND3_X1  g127(.A1(new_n297), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g128(.A1(new_n252), .A2(new_n253), .A3(new_n313), .ZN(new_n329));
  OAI21_X1  g129(.A(new_n329), .B1(new_n255), .B2(new_n313), .ZN(new_n330));
  INV_X1    g130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g131(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g132(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g134(.A1(new_n334), .A2(G33), .ZN(new_n335));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g136(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n337));
  OAI211_X1 g137(.A(KEYINPUT7), .B(new_n207), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n339));
  AND2_X1   g139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n335), .ZN(new_n341));
  AOI21_X1  g141(.A(KEYINPUT7), .B1(new_n341), .B2(new_n207), .ZN(new_n342));
  INV_X1    g142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g143(.A(new_n343), .B1(new_n338), .B2(new_n339), .ZN(new_n344));
  OAI21_X1  g144(.A(G68), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  OR2_X1    g145(.A1(new_n345), .A2(KEYINPUT80), .ZN(new_n346));
  INV_X1    g146(.A(G68), .ZN(new_n347));
  NOR2_X1   g147(.A1(new_n218), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g148(.A(G20), .B1(new_n348), .B2(new_n201), .ZN(new_n349));
  INV_X1    g149(.A(G159), .ZN(new_n350));
  OAI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n258), .ZN(new_n351));
  AOI21_X1  g151(.A(new_n351), .B1(new_n345), .B2(KEYINPUT80), .ZN(new_n352));
  AOI21_X1  g152(.A(KEYINPUT16), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g153(.A(new_n351), .B(KEYINPUT77), .ZN(new_n354));
  AND3_X1   g154(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n355));
  OAI21_X1  g155(.A(G68), .B1(new_n355), .B2(new_n342), .ZN(new_n356));
  AND2_X1   g156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g157(.A1(new_n357), .A2(KEYINPUT16), .ZN(new_n358));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n251), .ZN(new_n359));
  OAI21_X1  g159(.A(new_n331), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g160(.A1(new_n286), .A2(new_n219), .ZN(new_n361));
  XOR2_X1   g161(.A(new_n361), .B(KEYINPUT81), .Z(new_n362));
  OR2_X1    g162(.A1(G223), .A2(G1698), .ZN(new_n363));
  OAI21_X1  g163(.A(new_n363), .B1(G226), .B2(new_n299), .ZN(new_n364));
  INV_X1    g164(.A(G87), .ZN(new_n365));
  OAI22_X1  g165(.A1(new_n364), .A2(new_n341), .B1(new_n257), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g166(.A(new_n284), .B1(new_n277), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g168(.A1(new_n368), .A2(G169), .ZN(new_n369));
  OAI21_X1  g169(.A(new_n369), .B1(new_n310), .B2(new_n368), .ZN(new_n370));
  NAND2_X1  g170(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g171(.A1(new_n371), .A2(KEYINPUT18), .ZN(new_n372));
  INV_X1    g172(.A(KEYINPUT18), .ZN(new_n373));
  NAND3_X1  g173(.A1(new_n360), .A2(new_n373), .A3(new_n370), .ZN(new_n374));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g175(.A1(new_n368), .A2(new_n291), .ZN(new_n376));
  AOI21_X1  g176(.A(new_n376), .B1(G200), .B2(new_n368), .ZN(new_n377));
  OAI211_X1 g177(.A(new_n377), .B(new_n331), .C1(new_n353), .C2(new_n359), .ZN(new_n378));
  XNOR2_X1  g178(.A(new_n378), .B(KEYINPUT17), .ZN(new_n379));
  INV_X1    g179(.A(new_n379), .ZN(new_n380));
  NOR3_X1   g180(.A1(new_n328), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g181(.A(new_n284), .B1(new_n287), .B2(G238), .ZN(new_n382));
  NAND4_X1  g182(.A1(new_n332), .A2(new_n335), .A3(G232), .A4(G1698), .ZN(new_n383));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g185(.A1(new_n270), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n386));
  NAND2_X1  g186(.A1(G33), .A2(G97), .ZN(new_n387));
  NAND3_X1  g187(.A1(new_n270), .A2(G226), .A3(new_n299), .ZN(new_n388));
  NAND4_X1  g188(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  AND3_X1   g189(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n277), .ZN(new_n390));
  AOI21_X1  g190(.A(KEYINPUT73), .B1(new_n389), .B2(new_n277), .ZN(new_n391));
  OAI21_X1  g191(.A(new_n382), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g192(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n393));
  INV_X1    g193(.A(KEYINPUT74), .ZN(new_n394));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n395));
  OAI211_X1 g195(.A(new_n382), .B(new_n395), .C1(new_n390), .C2(new_n391), .ZN(new_n396));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g197(.A1(new_n392), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g198(.A1(new_n397), .A2(G200), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g199(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n347), .ZN(new_n400));
  OAI21_X1  g200(.A(new_n400), .B1(new_n262), .B2(new_n272), .ZN(new_n401));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n402));
  OR3_X1    g202(.A1(new_n255), .A2(KEYINPUT12), .A3(G68), .ZN(new_n403));
  OAI21_X1  g203(.A(KEYINPUT12), .B1(new_n255), .B2(G68), .ZN(new_n404));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g205(.A(new_n252), .ZN(new_n406));
  NAND2_X1  g206(.A1(new_n253), .A2(G68), .ZN(new_n407));
  OAI211_X1 g207(.A(new_n402), .B(new_n405), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g208(.A(KEYINPUT11), .B1(new_n401), .B2(new_n251), .ZN(new_n409));
  OR2_X1    g209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g210(.A(new_n291), .B1(new_n392), .B2(KEYINPUT13), .ZN(new_n411));
  AOI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n396), .ZN(new_n412));
  NAND2_X1  g212(.A1(new_n399), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g213(.A1(new_n413), .A2(KEYINPUT75), .ZN(new_n414));
  NOR2_X1   g214(.A1(new_n413), .A2(KEYINPUT75), .ZN(new_n415));
  NOR2_X1   g215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g216(.A1(new_n393), .A2(G179), .A3(new_n396), .ZN(new_n417));
  INV_X1    g217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g218(.A1(new_n397), .A2(G169), .A3(new_n398), .ZN(new_n419));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n420));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g221(.A1(new_n397), .A2(KEYINPUT14), .A3(G169), .A4(new_n398), .ZN(new_n422));
  AOI21_X1  g222(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g223(.A(new_n423), .B(KEYINPUT76), .ZN(new_n424));
  AOI21_X1  g224(.A(new_n416), .B1(new_n424), .B2(new_n410), .ZN(new_n425));
  NAND2_X1  g225(.A1(new_n381), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g226(.A(new_n252), .B1(G1), .B2(new_n257), .ZN(new_n427));
  AOI21_X1  g227(.A(KEYINPUT25), .B1(new_n249), .B2(new_n220), .ZN(new_n428));
  NAND3_X1  g228(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n429));
  INV_X1    g229(.A(new_n429), .ZN(new_n430));
  OAI22_X1  g230(.A1(new_n427), .A2(new_n220), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g231(.A(KEYINPUT22), .ZN(new_n432));
  NAND2_X1  g232(.A1(new_n270), .A2(new_n207), .ZN(new_n433));
  OAI211_X1 g233(.A(KEYINPUT87), .B(new_n432), .C1(new_n433), .C2(new_n365), .ZN(new_n434));
  XOR2_X1   g234(.A(KEYINPUT89), .B(KEYINPUT23), .Z(new_n435));
  OAI21_X1  g235(.A(new_n435), .B1(new_n207), .B2(new_n301), .ZN(new_n436));
  NOR3_X1   g236(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n437));
  NAND2_X1  g237(.A1(G33), .A2(G116), .ZN(new_n438));
  OR3_X1    g238(.A1(new_n438), .A2(KEYINPUT88), .A3(G20), .ZN(new_n439));
  OAI21_X1  g239(.A(KEYINPUT88), .B1(new_n438), .B2(G20), .ZN(new_n440));
  AOI21_X1  g240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g241(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n442));
  NAND4_X1  g242(.A1(new_n270), .A2(new_n442), .A3(new_n207), .A4(G87), .ZN(new_n443));
  NAND4_X1  g243(.A1(new_n434), .A2(new_n436), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  XNOR2_X1  g244(.A(new_n444), .B(KEYINPUT24), .ZN(new_n445));
  AOI21_X1  g245(.A(new_n431), .B1(new_n445), .B2(new_n251), .ZN(new_n446));
  INV_X1    g246(.A(new_n446), .ZN(new_n447));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n448));
  OAI211_X1 g248(.A(new_n206), .B(G45), .C1(new_n448), .C2(G41), .ZN(new_n449));
  INV_X1    g249(.A(new_n280), .ZN(new_n450));
  AOI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n448), .ZN(new_n451));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n277), .ZN(new_n452));
  NAND3_X1  g252(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n453));
  INV_X1    g253(.A(G294), .ZN(new_n454));
  INV_X1    g254(.A(G250), .ZN(new_n455));
  OAI221_X1 g255(.A(new_n453), .B1(new_n257), .B2(new_n454), .C1(new_n300), .C2(new_n455), .ZN(new_n456));
  AOI22_X1  g256(.A1(G264), .A2(new_n452), .B1(new_n456), .B2(new_n277), .ZN(new_n457));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n279), .ZN(new_n458));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g259(.A1(new_n459), .A2(G200), .ZN(new_n460));
  OAI21_X1  g260(.A(new_n460), .B1(new_n291), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n461), .ZN(new_n462));
  INV_X1    g262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g263(.A1(new_n341), .A2(G1698), .ZN(new_n464));
  NAND3_X1  g264(.A1(new_n464), .A2(KEYINPUT4), .A3(G244), .ZN(new_n465));
  NAND2_X1  g265(.A1(G33), .A2(G283), .ZN(new_n466));
  OAI211_X1 g266(.A(new_n465), .B(new_n466), .C1(new_n455), .C2(new_n304), .ZN(new_n467));
  AOI21_X1  g267(.A(KEYINPUT4), .B1(new_n464), .B2(G244), .ZN(new_n468));
  OAI21_X1  g268(.A(new_n277), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g269(.A1(new_n452), .A2(G257), .B1(new_n279), .B2(new_n451), .ZN(new_n470));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  OAI21_X1  g272(.A(new_n472), .B1(new_n291), .B2(new_n471), .ZN(new_n473));
  MUX2_X1   g273(.A(new_n255), .B(new_n427), .S(G97), .Z(new_n474));
  OAI21_X1  g274(.A(new_n301), .B1(new_n340), .B2(new_n344), .ZN(new_n475));
  NAND3_X1  g275(.A1(new_n220), .A2(KEYINPUT6), .A3(G97), .ZN(new_n476));
  XOR2_X1   g276(.A(G97), .B(G107), .Z(new_n477));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n479));
  AND2_X1   g279(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g280(.A(new_n474), .B1(new_n480), .B2(new_n312), .ZN(new_n481));
  OR2_X1    g281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g282(.A1(new_n427), .A2(new_n365), .ZN(new_n483));
  XNOR2_X1  g283(.A(new_n483), .B(KEYINPUT82), .ZN(new_n484));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n485));
  INV_X1    g285(.A(G97), .ZN(new_n486));
  OAI21_X1  g286(.A(new_n485), .B1(new_n262), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g287(.A1(new_n302), .A2(new_n365), .A3(new_n486), .ZN(new_n488));
  OAI21_X1  g288(.A(new_n207), .B1(new_n387), .B2(new_n485), .ZN(new_n489));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g290(.A(new_n487), .B(new_n490), .C1(new_n347), .C2(new_n433), .ZN(new_n491));
  AOI22_X1  g291(.A1(new_n491), .A2(new_n251), .B1(new_n249), .B2(new_n315), .ZN(new_n492));
  NAND2_X1  g292(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  INV_X1    g293(.A(G244), .ZN(new_n494));
  OAI221_X1 g294(.A(new_n438), .B1(new_n304), .B2(new_n494), .C1(new_n305), .C2(new_n300), .ZN(new_n495));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n277), .ZN(new_n496));
  NAND2_X1  g296(.A1(new_n206), .A2(G45), .ZN(new_n497));
  AOI21_X1  g297(.A(new_n277), .B1(new_n455), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g298(.A(new_n498), .B1(G274), .B2(new_n497), .ZN(new_n499));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g301(.A(new_n493), .B1(G190), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g302(.A1(new_n500), .A2(G200), .ZN(new_n503));
  NOR2_X1   g303(.A1(new_n500), .A2(G179), .ZN(new_n504));
  AOI21_X1  g304(.A(new_n504), .B1(new_n294), .B2(new_n500), .ZN(new_n505));
  OAI21_X1  g305(.A(new_n492), .B1(new_n315), .B2(new_n427), .ZN(new_n506));
  AOI22_X1  g306(.A1(new_n502), .A2(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g307(.A1(new_n471), .A2(G179), .ZN(new_n508));
  AOI21_X1  g308(.A(new_n508), .B1(new_n294), .B2(new_n471), .ZN(new_n509));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n481), .ZN(new_n510));
  NAND4_X1  g310(.A1(new_n463), .A2(new_n482), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g311(.A1(new_n459), .A2(new_n294), .ZN(new_n512));
  OAI21_X1  g312(.A(new_n512), .B1(G179), .B2(new_n459), .ZN(new_n513));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n446), .ZN(new_n514));
  INV_X1    g314(.A(new_n514), .ZN(new_n515));
  MUX2_X1   g315(.A(new_n255), .B(new_n427), .S(G116), .Z(new_n516));
  NOR2_X1   g316(.A1(new_n207), .A2(G116), .ZN(new_n517));
  OAI21_X1  g317(.A(KEYINPUT84), .B1(new_n312), .B2(new_n517), .ZN(new_n518));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n519));
  OAI211_X1 g319(.A(new_n251), .B(new_n519), .C1(new_n207), .C2(G116), .ZN(new_n520));
  OAI211_X1 g320(.A(new_n466), .B(new_n207), .C1(G33), .C2(new_n486), .ZN(new_n521));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OR2_X1    g322(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n523));
  NAND2_X1  g323(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n524));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g325(.A(new_n516), .B(new_n525), .C1(new_n523), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g326(.A1(new_n452), .A2(G270), .ZN(new_n527));
  NAND3_X1  g327(.A1(new_n270), .A2(G257), .A3(new_n299), .ZN(new_n528));
  XNOR2_X1  g328(.A(KEYINPUT83), .B(G303), .ZN(new_n529));
  OAI221_X1 g329(.A(new_n528), .B1(new_n270), .B2(new_n529), .C1(new_n304), .C2(new_n221), .ZN(new_n530));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n277), .ZN(new_n531));
  NAND3_X1  g331(.A1(new_n527), .A2(new_n531), .A3(new_n458), .ZN(new_n532));
  AND3_X1   g332(.A1(new_n526), .A2(G169), .A3(new_n532), .ZN(new_n533));
  INV_X1    g333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g334(.A1(new_n534), .A2(KEYINPUT86), .ZN(new_n535));
  OR2_X1    g335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g336(.A1(new_n532), .A2(new_n310), .ZN(new_n537));
  AOI22_X1  g337(.A1(new_n533), .A2(new_n535), .B1(new_n526), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g338(.A1(new_n532), .A2(G200), .ZN(new_n539));
  OAI21_X1  g339(.A(new_n539), .B1(new_n291), .B2(new_n532), .ZN(new_n540));
  OR2_X1    g340(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  NAND4_X1  g341(.A1(new_n515), .A2(new_n536), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  NOR3_X1   g342(.A1(new_n426), .A2(new_n511), .A3(new_n542), .ZN(G372));
  OR2_X1    g343(.A1(new_n414), .A2(new_n415), .ZN(new_n544));
  INV_X1    g344(.A(new_n323), .ZN(new_n545));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g346(.A1(new_n421), .A2(new_n422), .ZN(new_n547));
  AOI21_X1  g347(.A(KEYINPUT76), .B1(new_n547), .B2(new_n417), .ZN(new_n548));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n549));
  AOI211_X1 g349(.A(new_n549), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n550));
  OAI21_X1  g350(.A(new_n410), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g351(.A(new_n380), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n553));
  INV_X1    g353(.A(new_n374), .ZN(new_n554));
  AOI21_X1  g354(.A(new_n373), .B1(new_n360), .B2(new_n370), .ZN(new_n555));
  OAI21_X1  g355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g356(.A1(new_n372), .A2(KEYINPUT90), .A3(new_n374), .ZN(new_n557));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g358(.A(new_n293), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n296), .ZN(new_n560));
  NAND2_X1  g360(.A1(new_n560), .A2(KEYINPUT91), .ZN(new_n561));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n562));
  NAND3_X1  g362(.A1(new_n559), .A2(new_n562), .A3(new_n296), .ZN(new_n563));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g364(.A(new_n426), .ZN(new_n565));
  INV_X1    g365(.A(new_n510), .ZN(new_n566));
  AND3_X1   g366(.A1(new_n566), .A2(KEYINPUT26), .A3(new_n507), .ZN(new_n567));
  AOI21_X1  g367(.A(KEYINPUT26), .B1(new_n566), .B2(new_n507), .ZN(new_n568));
  NOR2_X1   g368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g369(.A1(new_n505), .A2(new_n506), .ZN(new_n570));
  NAND2_X1  g370(.A1(new_n536), .A2(new_n538), .ZN(new_n571));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n514), .ZN(new_n572));
  OAI21_X1  g372(.A(new_n570), .B1(new_n511), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g373(.A(new_n565), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g374(.A1(new_n564), .A2(new_n574), .ZN(G369));
  NAND3_X1  g375(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n576));
  XNOR2_X1  g376(.A(new_n576), .B(KEYINPUT92), .ZN(new_n577));
  INV_X1    g377(.A(new_n577), .ZN(new_n578));
  OR2_X1    g378(.A1(new_n578), .A2(KEYINPUT27), .ZN(new_n579));
  NAND2_X1  g379(.A1(new_n578), .A2(KEYINPUT27), .ZN(new_n580));
  NAND3_X1  g380(.A1(new_n579), .A2(G213), .A3(new_n580), .ZN(new_n581));
  INV_X1    g381(.A(G343), .ZN(new_n582));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n526), .ZN(new_n584));
  XOR2_X1   g384(.A(new_n584), .B(KEYINPUT93), .Z(new_n585));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g386(.A(new_n586), .B(KEYINPUT94), .ZN(new_n587));
  INV_X1    g387(.A(new_n585), .ZN(new_n588));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n541), .ZN(new_n589));
  OAI21_X1  g389(.A(new_n587), .B1(new_n571), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g390(.A1(new_n590), .A2(G330), .ZN(new_n591));
  INV_X1    g391(.A(new_n591), .ZN(new_n592));
  INV_X1    g392(.A(new_n583), .ZN(new_n593));
  NAND2_X1  g393(.A1(new_n514), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g394(.A1(new_n446), .A2(new_n593), .ZN(new_n595));
  NOR2_X1   g395(.A1(new_n462), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g396(.A(new_n594), .B1(new_n596), .B2(new_n514), .ZN(new_n597));
  XNOR2_X1  g397(.A(new_n597), .B(KEYINPUT95), .ZN(new_n598));
  NAND2_X1  g398(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g399(.A1(new_n571), .A2(new_n593), .ZN(new_n600));
  XOR2_X1   g400(.A(new_n600), .B(KEYINPUT96), .Z(new_n601));
  AOI22_X1  g401(.A1(new_n598), .A2(new_n601), .B1(new_n514), .B2(new_n593), .ZN(new_n602));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n602), .ZN(G399));
  NOR2_X1   g403(.A1(new_n488), .A2(G116), .ZN(new_n604));
  NAND2_X1  g404(.A1(new_n210), .A2(new_n280), .ZN(new_n605));
  NAND3_X1  g405(.A1(new_n604), .A2(G1), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g406(.A(new_n606), .B1(new_n216), .B2(new_n605), .ZN(new_n607));
  XNOR2_X1  g407(.A(new_n607), .B(KEYINPUT28), .ZN(new_n608));
  OAI21_X1  g408(.A(new_n593), .B1(new_n569), .B2(new_n573), .ZN(new_n609));
  XOR2_X1   g409(.A(new_n609), .B(KEYINPUT29), .Z(new_n610));
  NOR3_X1   g410(.A1(new_n511), .A2(new_n542), .A3(new_n583), .ZN(new_n611));
  INV_X1    g411(.A(new_n611), .ZN(new_n612));
  INV_X1    g412(.A(KEYINPUT30), .ZN(new_n613));
  NAND3_X1  g413(.A1(new_n537), .A2(new_n457), .A3(new_n501), .ZN(new_n614));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n471), .ZN(new_n615));
  AND2_X1   g415(.A1(new_n532), .A2(new_n310), .ZN(new_n616));
  NAND4_X1  g416(.A1(new_n616), .A2(new_n471), .A3(new_n459), .A4(new_n500), .ZN(new_n617));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g418(.A1(new_n614), .A2(new_n613), .A3(new_n471), .ZN(new_n619));
  OAI21_X1  g419(.A(new_n583), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g420(.A(new_n620), .B(KEYINPUT31), .ZN(new_n621));
  NAND2_X1  g421(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g422(.A1(new_n622), .A2(G330), .ZN(new_n623));
  NAND2_X1  g423(.A1(new_n610), .A2(new_n623), .ZN(new_n624));
  INV_X1    g424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g425(.A(new_n608), .B1(new_n625), .B2(G1), .ZN(G364));
  INV_X1    g426(.A(new_n605), .ZN(new_n627));
  NOR2_X1   g427(.A1(new_n248), .A2(G20), .ZN(new_n628));
  AOI21_X1  g428(.A(new_n206), .B1(new_n628), .B2(G45), .ZN(new_n629));
  INV_X1    g429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g431(.A1(new_n592), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g432(.A1(new_n590), .A2(G330), .ZN(new_n633));
  INV_X1    g433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g434(.A1(G13), .A2(G33), .ZN(new_n635));
  INV_X1    g435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  INV_X1    g437(.A(new_n637), .ZN(new_n638));
  OR2_X1    g438(.A1(new_n590), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g439(.A1(new_n210), .A2(new_n270), .ZN(new_n640));
  INV_X1    g440(.A(G355), .ZN(new_n641));
  OAI22_X1  g441(.A1(new_n640), .A2(new_n641), .B1(G116), .B2(new_n210), .ZN(new_n642));
  OR2_X1    g442(.A1(new_n243), .A2(new_n281), .ZN(new_n643));
  NAND2_X1  g443(.A1(new_n210), .A2(new_n341), .ZN(new_n644));
  INV_X1    g444(.A(new_n216), .ZN(new_n645));
  AOI21_X1  g445(.A(new_n644), .B1(new_n281), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g446(.A(new_n642), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g447(.A1(new_n294), .A2(KEYINPUT97), .ZN(new_n648));
  INV_X1    g448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g449(.A(new_n207), .B1(KEYINPUT97), .B2(new_n294), .ZN(new_n650));
  AOI21_X1  g450(.A(new_n213), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n637), .ZN(new_n652));
  INV_X1    g452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g453(.A(new_n631), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g454(.A1(new_n207), .A2(G179), .ZN(new_n655));
  NAND3_X1  g455(.A1(new_n655), .A2(G190), .A3(G200), .ZN(new_n656));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n365), .ZN(new_n657));
  NOR2_X1   g457(.A1(G190), .A2(G200), .ZN(new_n658));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g460(.A1(new_n660), .A2(G159), .ZN(new_n661));
  NOR2_X1   g461(.A1(new_n661), .A2(KEYINPUT32), .ZN(new_n662));
  NOR2_X1   g462(.A1(new_n207), .A2(new_n310), .ZN(new_n663));
  NAND2_X1  g463(.A1(new_n663), .A2(G200), .ZN(new_n664));
  NOR2_X1   g464(.A1(new_n664), .A2(G190), .ZN(new_n665));
  AOI211_X1 g465(.A(new_n657), .B(new_n662), .C1(G68), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n658), .ZN(new_n667));
  OAI21_X1  g467(.A(new_n270), .B1(new_n667), .B2(new_n272), .ZN(new_n668));
  NAND3_X1  g468(.A1(new_n663), .A2(G190), .A3(new_n324), .ZN(new_n669));
  INV_X1    g469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g470(.A(new_n668), .B1(G58), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n291), .A3(G200), .ZN(new_n672));
  INV_X1    g472(.A(new_n672), .ZN(new_n673));
  AOI22_X1  g473(.A1(new_n661), .A2(KEYINPUT32), .B1(G107), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g474(.A1(new_n291), .A2(G179), .A3(G200), .ZN(new_n675));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n207), .ZN(new_n676));
  INV_X1    g476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g477(.A1(new_n664), .A2(new_n291), .ZN(new_n678));
  AOI22_X1  g478(.A1(G97), .A2(new_n677), .B1(new_n678), .B2(G50), .ZN(new_n679));
  NAND4_X1  g479(.A1(new_n666), .A2(new_n671), .A3(new_n674), .A4(new_n679), .ZN(new_n680));
  INV_X1    g480(.A(G322), .ZN(new_n681));
  NOR2_X1   g481(.A1(new_n669), .A2(new_n681), .ZN(new_n682));
  INV_X1    g482(.A(G311), .ZN(new_n683));
  OAI21_X1  g483(.A(new_n341), .B1(new_n667), .B2(new_n683), .ZN(new_n684));
  AOI211_X1 g484(.A(new_n682), .B(new_n684), .C1(G329), .C2(new_n660), .ZN(new_n685));
  NAND2_X1  g485(.A1(new_n678), .A2(G326), .ZN(new_n686));
  XNOR2_X1  g486(.A(KEYINPUT33), .B(G317), .ZN(new_n687));
  INV_X1    g487(.A(new_n656), .ZN(new_n688));
  AOI22_X1  g488(.A1(new_n665), .A2(new_n687), .B1(new_n688), .B2(G303), .ZN(new_n689));
  AOI22_X1  g489(.A1(new_n677), .A2(G294), .B1(new_n673), .B2(G283), .ZN(new_n690));
  NAND4_X1  g490(.A1(new_n685), .A2(new_n686), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g491(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g492(.A(new_n654), .B1(new_n692), .B2(new_n651), .ZN(new_n693));
  AOI22_X1  g493(.A1(new_n632), .A2(new_n634), .B1(new_n639), .B2(new_n693), .ZN(new_n694));
  INV_X1    g494(.A(new_n694), .ZN(G396));
  NOR2_X1   g495(.A1(new_n323), .A2(new_n583), .ZN(new_n696));
  OAI21_X1  g496(.A(new_n327), .B1(new_n320), .B2(new_n593), .ZN(new_n697));
  AOI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n323), .ZN(new_n698));
  INV_X1    g498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g499(.A1(new_n609), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g500(.A(new_n593), .B(new_n698), .C1(new_n569), .C2(new_n573), .ZN(new_n701));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g502(.A(new_n631), .B1(new_n702), .B2(new_n623), .ZN(new_n703));
  OAI21_X1  g503(.A(new_n703), .B1(new_n623), .B2(new_n702), .ZN(new_n704));
  INV_X1    g504(.A(new_n631), .ZN(new_n705));
  NOR2_X1   g505(.A1(new_n651), .A2(new_n635), .ZN(new_n706));
  XOR2_X1   g506(.A(new_n706), .B(KEYINPUT98), .Z(new_n707));
  INV_X1    g507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n272), .ZN(new_n709));
  INV_X1    g509(.A(new_n651), .ZN(new_n710));
  AOI22_X1  g510(.A1(new_n670), .A2(G294), .B1(new_n660), .B2(G311), .ZN(new_n711));
  INV_X1    g511(.A(G116), .ZN(new_n712));
  OAI211_X1 g512(.A(new_n711), .B(new_n341), .C1(new_n712), .C2(new_n667), .ZN(new_n713));
  AOI22_X1  g513(.A1(new_n678), .A2(G303), .B1(new_n673), .B2(G87), .ZN(new_n714));
  OAI21_X1  g514(.A(new_n714), .B1(new_n220), .B2(new_n656), .ZN(new_n715));
  INV_X1    g515(.A(new_n665), .ZN(new_n716));
  INV_X1    g516(.A(G283), .ZN(new_n717));
  OAI22_X1  g517(.A1(new_n716), .A2(new_n717), .B1(new_n486), .B2(new_n676), .ZN(new_n718));
  NOR3_X1   g518(.A1(new_n713), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g519(.A1(new_n672), .A2(new_n347), .ZN(new_n720));
  INV_X1    g520(.A(G132), .ZN(new_n721));
  OAI221_X1 g521(.A(new_n270), .B1(new_n659), .B2(new_n721), .C1(new_n202), .C2(new_n656), .ZN(new_n722));
  AOI211_X1 g522(.A(new_n720), .B(new_n722), .C1(G58), .C2(new_n677), .ZN(new_n723));
  XNOR2_X1  g523(.A(new_n723), .B(KEYINPUT99), .ZN(new_n724));
  INV_X1    g524(.A(new_n667), .ZN(new_n725));
  AOI22_X1  g525(.A1(new_n670), .A2(G143), .B1(new_n725), .B2(G159), .ZN(new_n726));
  INV_X1    g526(.A(G150), .ZN(new_n727));
  INV_X1    g527(.A(G137), .ZN(new_n728));
  INV_X1    g528(.A(new_n678), .ZN(new_n729));
  OAI221_X1 g529(.A(new_n726), .B1(new_n716), .B2(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g530(.A(new_n730), .B(KEYINPUT34), .ZN(new_n731));
  AOI21_X1  g531(.A(new_n719), .B1(new_n724), .B2(new_n731), .ZN(new_n732));
  OAI221_X1 g532(.A(new_n709), .B1(new_n710), .B2(new_n732), .C1(new_n698), .C2(new_n636), .ZN(new_n733));
  AND2_X1   g533(.A1(new_n704), .A2(new_n733), .ZN(new_n734));
  INV_X1    g534(.A(new_n734), .ZN(G384));
  AOI211_X1 g535(.A(new_n712), .B(new_n215), .C1(new_n478), .C2(KEYINPUT35), .ZN(new_n736));
  OAI21_X1  g536(.A(new_n736), .B1(KEYINPUT35), .B2(new_n478), .ZN(new_n737));
  XNOR2_X1  g537(.A(new_n737), .B(KEYINPUT36), .ZN(new_n738));
  OAI21_X1  g538(.A(G77), .B1(new_n218), .B2(new_n347), .ZN(new_n739));
  OAI22_X1  g539(.A1(new_n739), .A2(new_n216), .B1(G50), .B2(new_n347), .ZN(new_n740));
  NAND3_X1  g540(.A1(new_n740), .A2(G1), .A3(new_n248), .ZN(new_n741));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g542(.A(new_n742), .B(KEYINPUT100), .Z(new_n743));
  INV_X1    g543(.A(KEYINPUT40), .ZN(new_n744));
  NOR2_X1   g544(.A1(new_n357), .A2(KEYINPUT16), .ZN(new_n745));
  OAI21_X1  g545(.A(new_n331), .B1(new_n359), .B2(new_n745), .ZN(new_n746));
  INV_X1    g546(.A(new_n581), .ZN(new_n747));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g548(.A1(new_n554), .A2(new_n555), .ZN(new_n749));
  AOI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n379), .ZN(new_n750));
  INV_X1    g550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g551(.A1(new_n360), .A2(new_n747), .ZN(new_n752));
  INV_X1    g552(.A(KEYINPUT37), .ZN(new_n753));
  NAND4_X1  g553(.A1(new_n371), .A2(new_n752), .A3(new_n753), .A4(new_n378), .ZN(new_n754));
  OAI21_X1  g554(.A(new_n746), .B1(new_n370), .B2(new_n747), .ZN(new_n755));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n378), .ZN(new_n756));
  NAND2_X1  g556(.A1(new_n756), .A2(KEYINPUT37), .ZN(new_n757));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g558(.A1(new_n751), .A2(KEYINPUT38), .A3(new_n758), .ZN(new_n759));
  INV_X1    g559(.A(KEYINPUT38), .ZN(new_n760));
  INV_X1    g560(.A(new_n758), .ZN(new_n761));
  OAI21_X1  g561(.A(new_n760), .B1(new_n750), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g563(.A(KEYINPUT31), .ZN(new_n764));
  XNOR2_X1  g564(.A(new_n620), .B(new_n764), .ZN(new_n765));
  OAI21_X1  g565(.A(new_n698), .B1(new_n765), .B2(new_n611), .ZN(new_n766));
  OAI211_X1 g566(.A(new_n410), .B(new_n583), .C1(new_n424), .C2(new_n416), .ZN(new_n767));
  NAND2_X1  g567(.A1(new_n410), .A2(new_n583), .ZN(new_n768));
  NAND3_X1  g568(.A1(new_n551), .A2(new_n544), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g569(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g570(.A(KEYINPUT102), .ZN(new_n771));
  OAI21_X1  g571(.A(new_n763), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g572(.A(KEYINPUT102), .B(new_n766), .C1(new_n767), .C2(new_n769), .ZN(new_n773));
  OAI21_X1  g573(.A(new_n744), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g574(.A1(new_n774), .A2(KEYINPUT103), .ZN(new_n775));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n776));
  OAI211_X1 g576(.A(new_n776), .B(new_n744), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g578(.A(new_n699), .B1(new_n612), .B2(new_n621), .ZN(new_n779));
  AND3_X1   g579(.A1(new_n551), .A2(new_n544), .A3(new_n768), .ZN(new_n780));
  AOI21_X1  g580(.A(new_n768), .B1(new_n551), .B2(new_n544), .ZN(new_n781));
  OAI21_X1  g581(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g582(.A(new_n752), .ZN(new_n783));
  OAI21_X1  g583(.A(new_n783), .B1(new_n558), .B2(new_n380), .ZN(new_n784));
  NAND3_X1  g584(.A1(new_n371), .A2(new_n752), .A3(new_n378), .ZN(new_n785));
  NAND2_X1  g585(.A1(new_n785), .A2(KEYINPUT37), .ZN(new_n786));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n754), .ZN(new_n787));
  AOI21_X1  g587(.A(KEYINPUT38), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g588(.A1(new_n750), .A2(new_n761), .A3(new_n760), .ZN(new_n789));
  OAI21_X1  g589(.A(KEYINPUT40), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g590(.A(new_n778), .B1(new_n782), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g591(.A1(new_n565), .A2(new_n622), .ZN(new_n792));
  AND2_X1   g592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  INV_X1    g594(.A(G330), .ZN(new_n795));
  NOR3_X1   g595(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g596(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g597(.A1(new_n424), .A2(new_n410), .A3(new_n593), .ZN(new_n798));
  XOR2_X1   g598(.A(new_n798), .B(KEYINPUT101), .Z(new_n799));
  NAND3_X1  g599(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT39), .ZN(new_n800));
  NOR2_X1   g600(.A1(new_n788), .A2(new_n789), .ZN(new_n801));
  OAI211_X1 g601(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(KEYINPUT39), .ZN(new_n802));
  NAND2_X1  g602(.A1(new_n767), .A2(new_n769), .ZN(new_n803));
  INV_X1    g603(.A(new_n696), .ZN(new_n804));
  NAND2_X1  g604(.A1(new_n701), .A2(new_n804), .ZN(new_n805));
  AND2_X1   g605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n763), .ZN(new_n807));
  NAND2_X1  g607(.A1(new_n558), .A2(new_n581), .ZN(new_n808));
  NAND3_X1  g608(.A1(new_n802), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g609(.A(new_n809), .ZN(new_n810));
  OR2_X1    g610(.A1(new_n610), .A2(new_n426), .ZN(new_n811));
  AND2_X1   g611(.A1(new_n564), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g612(.A(new_n810), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n813), .ZN(new_n814));
  INV_X1    g614(.A(new_n813), .ZN(new_n815));
  OAI22_X1  g615(.A1(new_n796), .A2(new_n815), .B1(new_n206), .B2(new_n628), .ZN(new_n816));
  OAI21_X1  g616(.A(new_n743), .B1(new_n814), .B2(new_n816), .ZN(G367));
  NAND2_X1  g617(.A1(new_n598), .A2(new_n601), .ZN(new_n818));
  NAND2_X1  g618(.A1(new_n566), .A2(new_n583), .ZN(new_n819));
  NAND2_X1  g619(.A1(new_n481), .A2(new_n583), .ZN(new_n820));
  NAND3_X1  g620(.A1(new_n482), .A2(new_n510), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g623(.A(KEYINPUT42), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g624(.A1(new_n821), .A2(new_n515), .ZN(new_n825));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n566), .ZN(new_n826));
  AOI21_X1  g626(.A(new_n583), .B1(new_n826), .B2(KEYINPUT105), .ZN(new_n827));
  OAI21_X1  g627(.A(new_n827), .B1(KEYINPUT105), .B2(new_n826), .ZN(new_n828));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g629(.A1(new_n829), .A2(KEYINPUT106), .ZN(new_n830));
  NOR3_X1   g630(.A1(new_n818), .A2(KEYINPUT42), .A3(new_n823), .ZN(new_n831));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g632(.A1(new_n829), .A2(KEYINPUT106), .ZN(new_n833));
  NAND2_X1  g633(.A1(new_n493), .A2(new_n583), .ZN(new_n834));
  NAND2_X1  g634(.A1(new_n507), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g635(.A(new_n835), .B1(new_n570), .B2(new_n834), .ZN(new_n836));
  AND2_X1   g636(.A1(new_n836), .A2(KEYINPUT104), .ZN(new_n837));
  NOR2_X1   g637(.A1(new_n836), .A2(KEYINPUT104), .ZN(new_n838));
  NOR3_X1   g638(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT43), .ZN(new_n839));
  NAND3_X1  g639(.A1(new_n832), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  INV_X1    g640(.A(KEYINPUT107), .ZN(new_n841));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g642(.A1(new_n832), .A2(KEYINPUT107), .A3(new_n833), .A4(new_n839), .ZN(new_n843));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g644(.A1(new_n832), .A2(new_n833), .ZN(new_n845));
  AOI21_X1  g645(.A(new_n839), .B1(KEYINPUT43), .B2(new_n836), .ZN(new_n846));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g648(.A1(new_n599), .A2(new_n823), .ZN(new_n849));
  INV_X1    g649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g650(.A1(new_n848), .A2(KEYINPUT108), .A3(new_n850), .ZN(new_n851));
  INV_X1    g651(.A(KEYINPUT108), .ZN(new_n852));
  AOI22_X1  g652(.A1(new_n842), .A2(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  OAI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n849), .ZN(new_n854));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n849), .ZN(new_n855));
  INV_X1    g655(.A(KEYINPUT45), .ZN(new_n856));
  INV_X1    g656(.A(new_n602), .ZN(new_n857));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n823), .ZN(new_n858));
  NAND3_X1  g658(.A1(new_n602), .A2(KEYINPUT45), .A3(new_n822), .ZN(new_n859));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g660(.A1(new_n857), .A2(KEYINPUT44), .A3(new_n823), .ZN(new_n861));
  INV_X1    g661(.A(KEYINPUT44), .ZN(new_n862));
  OAI21_X1  g662(.A(new_n862), .B1(new_n602), .B2(new_n822), .ZN(new_n863));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n599), .A3(new_n864), .ZN(new_n865));
  INV_X1    g665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g666(.A(new_n599), .B1(new_n860), .B2(new_n864), .ZN(new_n867));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g668(.A1(new_n598), .A2(new_n601), .ZN(new_n869));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n818), .ZN(new_n870));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n591), .ZN(new_n871));
  NAND3_X1  g671(.A1(new_n592), .A2(new_n818), .A3(new_n869), .ZN(new_n872));
  NAND4_X1  g672(.A1(new_n871), .A2(new_n610), .A3(new_n872), .A4(new_n623), .ZN(new_n873));
  INV_X1    g673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g674(.A(new_n624), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g675(.A(new_n605), .B(KEYINPUT41), .ZN(new_n876));
  OAI21_X1  g676(.A(new_n629), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g677(.A1(new_n851), .A2(new_n854), .A3(new_n855), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g678(.A1(new_n235), .A2(new_n644), .ZN(new_n879));
  OAI21_X1  g679(.A(new_n652), .B1(new_n210), .B2(new_n315), .ZN(new_n880));
  OAI21_X1  g680(.A(new_n631), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI22_X1  g681(.A1(new_n716), .A2(new_n350), .B1(new_n672), .B2(new_n272), .ZN(new_n882));
  AOI21_X1  g682(.A(new_n882), .B1(G58), .B2(new_n688), .ZN(new_n883));
  OAI22_X1  g683(.A1(new_n669), .A2(new_n727), .B1(new_n659), .B2(new_n728), .ZN(new_n884));
  AOI211_X1 g684(.A(new_n341), .B(new_n884), .C1(G50), .C2(new_n725), .ZN(new_n885));
  NAND2_X1  g685(.A1(new_n678), .A2(G143), .ZN(new_n886));
  NAND2_X1  g686(.A1(new_n677), .A2(G68), .ZN(new_n887));
  NAND4_X1  g687(.A1(new_n883), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g688(.A1(new_n656), .A2(new_n712), .ZN(new_n889));
  NOR2_X1   g689(.A1(new_n889), .A2(KEYINPUT46), .ZN(new_n890));
  XOR2_X1   g690(.A(new_n890), .B(KEYINPUT110), .Z(new_n891));
  NAND2_X1  g691(.A1(new_n673), .A2(G97), .ZN(new_n892));
  OAI21_X1  g692(.A(new_n892), .B1(new_n716), .B2(new_n454), .ZN(new_n893));
  AOI21_X1  g693(.A(new_n893), .B1(G311), .B2(new_n678), .ZN(new_n894));
  INV_X1    g694(.A(G317), .ZN(new_n895));
  OAI221_X1 g695(.A(new_n341), .B1(new_n659), .B2(new_n895), .C1(new_n669), .C2(new_n529), .ZN(new_n896));
  AOI21_X1  g696(.A(new_n896), .B1(KEYINPUT46), .B2(new_n889), .ZN(new_n897));
  NAND3_X1  g697(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  OAI22_X1  g698(.A1(new_n676), .A2(new_n302), .B1(new_n667), .B2(new_n717), .ZN(new_n899));
  XOR2_X1   g699(.A(new_n899), .B(KEYINPUT109), .Z(new_n900));
  OAI21_X1  g700(.A(new_n888), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g701(.A(new_n901), .B(KEYINPUT47), .ZN(new_n902));
  AOI21_X1  g702(.A(new_n881), .B1(new_n902), .B2(new_n651), .ZN(new_n903));
  OAI21_X1  g703(.A(new_n903), .B1(new_n836), .B2(new_n638), .ZN(new_n904));
  NAND2_X1  g704(.A1(new_n878), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g705(.A(new_n905), .B(KEYINPUT111), .Z(new_n906));
  INV_X1    g706(.A(new_n906), .ZN(G387));
  NAND2_X1  g707(.A1(new_n871), .A2(new_n872), .ZN(new_n908));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n624), .ZN(new_n909));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n873), .A3(new_n627), .ZN(new_n910));
  NAND3_X1  g710(.A1(new_n871), .A2(new_n872), .A3(new_n630), .ZN(new_n911));
  OAI22_X1  g711(.A1(new_n604), .A2(new_n640), .B1(G107), .B2(new_n210), .ZN(new_n912));
  NOR2_X1   g712(.A1(new_n239), .A2(new_n281), .ZN(new_n913));
  XNOR2_X1  g713(.A(new_n913), .B(KEYINPUT112), .ZN(new_n914));
  INV_X1    g714(.A(new_n604), .ZN(new_n915));
  AOI211_X1 g715(.A(G45), .B(new_n915), .C1(G68), .C2(G77), .ZN(new_n916));
  NOR2_X1   g716(.A1(new_n263), .A2(G50), .ZN(new_n917));
  XNOR2_X1  g717(.A(new_n917), .B(KEYINPUT50), .ZN(new_n918));
  AOI21_X1  g718(.A(new_n644), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g719(.A(new_n912), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g720(.A(new_n631), .B1(new_n920), .B2(new_n653), .ZN(new_n921));
  INV_X1    g721(.A(new_n315), .ZN(new_n922));
  AOI22_X1  g722(.A1(new_n922), .A2(new_n677), .B1(new_n665), .B2(new_n313), .ZN(new_n923));
  NAND2_X1  g723(.A1(new_n688), .A2(G77), .ZN(new_n924));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n892), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g725(.A1(new_n670), .A2(G50), .B1(new_n660), .B2(G150), .ZN(new_n926));
  OAI211_X1 g726(.A(new_n926), .B(new_n270), .C1(new_n347), .C2(new_n667), .ZN(new_n927));
  NOR3_X1   g727(.A1(new_n729), .A2(KEYINPUT113), .A3(new_n350), .ZN(new_n928));
  INV_X1    g728(.A(KEYINPUT113), .ZN(new_n929));
  AOI21_X1  g729(.A(new_n929), .B1(new_n678), .B2(G159), .ZN(new_n930));
  NOR4_X1   g730(.A1(new_n925), .A2(new_n927), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  XNOR2_X1  g731(.A(new_n931), .B(KEYINPUT114), .ZN(new_n932));
  INV_X1    g732(.A(new_n529), .ZN(new_n933));
  AOI22_X1  g733(.A1(new_n670), .A2(G317), .B1(new_n725), .B2(new_n933), .ZN(new_n934));
  OAI221_X1 g734(.A(new_n934), .B1(new_n716), .B2(new_n683), .C1(new_n681), .C2(new_n729), .ZN(new_n935));
  INV_X1    g735(.A(KEYINPUT48), .ZN(new_n936));
  OR2_X1    g736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  AOI22_X1  g738(.A1(new_n677), .A2(G283), .B1(new_n688), .B2(G294), .ZN(new_n939));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g740(.A(new_n940), .B(KEYINPUT115), .ZN(new_n941));
  NAND2_X1  g741(.A1(new_n941), .A2(KEYINPUT49), .ZN(new_n942));
  AOI21_X1  g742(.A(new_n270), .B1(new_n660), .B2(G326), .ZN(new_n943));
  OAI211_X1 g743(.A(new_n942), .B(new_n943), .C1(new_n712), .C2(new_n672), .ZN(new_n944));
  NOR2_X1   g744(.A1(new_n941), .A2(KEYINPUT49), .ZN(new_n945));
  OAI21_X1  g745(.A(new_n932), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g746(.A(new_n921), .B1(new_n946), .B2(new_n651), .ZN(new_n947));
  OAI21_X1  g747(.A(new_n947), .B1(new_n598), .B2(new_n638), .ZN(new_n948));
  AND2_X1   g748(.A1(new_n911), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g749(.A1(new_n910), .A2(new_n949), .ZN(G393));
  OAI21_X1  g750(.A(new_n873), .B1(new_n866), .B2(new_n867), .ZN(new_n951));
  INV_X1    g751(.A(new_n867), .ZN(new_n952));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n874), .A3(new_n865), .ZN(new_n953));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n953), .A3(new_n627), .ZN(new_n954));
  NOR2_X1   g754(.A1(new_n246), .A2(new_n644), .ZN(new_n955));
  OAI21_X1  g755(.A(new_n652), .B1(new_n486), .B2(new_n210), .ZN(new_n956));
  OAI21_X1  g756(.A(new_n631), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g757(.A1(new_n822), .A2(new_n638), .ZN(new_n958));
  AOI22_X1  g758(.A1(G150), .A2(new_n678), .B1(new_n670), .B2(G159), .ZN(new_n959));
  XNOR2_X1  g759(.A(new_n959), .B(KEYINPUT51), .ZN(new_n960));
  AOI21_X1  g760(.A(new_n341), .B1(new_n660), .B2(G143), .ZN(new_n961));
  OAI21_X1  g761(.A(new_n961), .B1(new_n263), .B2(new_n667), .ZN(new_n962));
  OAI22_X1  g762(.A1(new_n716), .A2(new_n202), .B1(new_n672), .B2(new_n365), .ZN(new_n963));
  OAI22_X1  g763(.A1(new_n676), .A2(new_n272), .B1(new_n656), .B2(new_n347), .ZN(new_n964));
  NOR4_X1   g764(.A1(new_n960), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g765(.A1(G317), .A2(new_n678), .B1(new_n670), .B2(G311), .ZN(new_n966));
  XNOR2_X1  g766(.A(new_n966), .B(KEYINPUT52), .ZN(new_n967));
  OAI221_X1 g767(.A(new_n341), .B1(new_n659), .B2(new_n681), .C1(new_n454), .C2(new_n667), .ZN(new_n968));
  OAI22_X1  g768(.A1(new_n220), .A2(new_n672), .B1(new_n656), .B2(new_n717), .ZN(new_n969));
  OAI22_X1  g769(.A1(new_n716), .A2(new_n529), .B1(new_n712), .B2(new_n676), .ZN(new_n970));
  NOR4_X1   g770(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g771(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  AOI211_X1 g772(.A(new_n957), .B(new_n958), .C1(new_n651), .C2(new_n972), .ZN(new_n973));
  AOI21_X1  g773(.A(new_n973), .B1(new_n868), .B2(new_n630), .ZN(new_n974));
  NAND2_X1  g774(.A1(new_n954), .A2(new_n974), .ZN(G390));
  XNOR2_X1  g775(.A(KEYINPUT54), .B(G143), .ZN(new_n976));
  OAI22_X1  g776(.A1(new_n669), .A2(new_n721), .B1(new_n667), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g777(.A(new_n341), .B(new_n977), .C1(G125), .C2(new_n660), .ZN(new_n978));
  NOR2_X1   g778(.A1(new_n656), .A2(new_n727), .ZN(new_n979));
  XNOR2_X1  g779(.A(new_n979), .B(KEYINPUT53), .ZN(new_n980));
  AOI22_X1  g780(.A1(new_n665), .A2(G137), .B1(new_n673), .B2(G50), .ZN(new_n981));
  NOR2_X1   g781(.A1(new_n676), .A2(new_n350), .ZN(new_n982));
  AOI21_X1  g782(.A(new_n982), .B1(G128), .B2(new_n678), .ZN(new_n983));
  NAND4_X1  g783(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g784(.A(new_n341), .B1(new_n669), .B2(new_n712), .ZN(new_n985));
  OAI22_X1  g785(.A1(new_n667), .A2(new_n486), .B1(new_n659), .B2(new_n454), .ZN(new_n986));
  NOR4_X1   g786(.A1(new_n985), .A2(new_n986), .A3(new_n657), .A4(new_n720), .ZN(new_n987));
  AOI22_X1  g787(.A1(G77), .A2(new_n677), .B1(new_n678), .B2(G283), .ZN(new_n988));
  OAI211_X1 g788(.A(new_n987), .B(new_n988), .C1(new_n302), .C2(new_n716), .ZN(new_n989));
  AOI21_X1  g789(.A(new_n710), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g790(.A(new_n705), .B(new_n990), .C1(new_n263), .C2(new_n708), .ZN(new_n991));
  XOR2_X1   g791(.A(new_n991), .B(KEYINPUT117), .Z(new_n992));
  OAI21_X1  g792(.A(new_n800), .B1(new_n801), .B2(KEYINPUT39), .ZN(new_n993));
  INV_X1    g793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n636), .ZN(new_n995));
  OAI21_X1  g795(.A(new_n993), .B1(new_n799), .B2(new_n806), .ZN(new_n996));
  OR3_X1    g796(.A1(new_n799), .A2(new_n801), .A3(new_n806), .ZN(new_n997));
  NAND3_X1  g797(.A1(new_n803), .A2(G330), .A3(new_n779), .ZN(new_n998));
  AND3_X1   g798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g799(.A(new_n998), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g802(.A(new_n995), .B1(new_n1002), .B2(new_n629), .ZN(new_n1003));
  OR2_X1    g803(.A1(new_n426), .A2(new_n623), .ZN(new_n1004));
  NAND2_X1  g804(.A1(new_n779), .A2(G330), .ZN(new_n1005));
  NAND3_X1  g805(.A1(new_n1005), .A2(new_n769), .A3(new_n767), .ZN(new_n1006));
  NAND2_X1  g806(.A1(new_n998), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n805), .ZN(new_n1008));
  NAND4_X1  g808(.A1(new_n998), .A2(new_n804), .A3(new_n1006), .A4(new_n701), .ZN(new_n1009));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g810(.A1(new_n812), .A2(KEYINPUT116), .A3(new_n1004), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g811(.A(KEYINPUT116), .ZN(new_n1012));
  INV_X1    g812(.A(new_n1010), .ZN(new_n1013));
  NAND3_X1  g813(.A1(new_n564), .A2(new_n811), .A3(new_n1004), .ZN(new_n1014));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g817(.A(new_n605), .B1(new_n1017), .B2(new_n1002), .ZN(new_n1018));
  NAND2_X1  g818(.A1(new_n1016), .A2(new_n1001), .ZN(new_n1019));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g820(.A(new_n1020), .ZN(G378));
  NOR2_X1   g821(.A1(new_n581), .A2(new_n265), .ZN(new_n1022));
  XNOR2_X1  g822(.A(new_n1022), .B(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g823(.A(new_n297), .B(new_n1023), .ZN(new_n1024));
  XOR2_X1   g824(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1025));
  XOR2_X1   g825(.A(new_n1024), .B(new_n1025), .Z(new_n1026));
  NAND2_X1  g826(.A1(new_n1026), .A2(new_n635), .ZN(new_n1027));
  OAI21_X1  g827(.A(new_n631), .B1(new_n707), .B2(G50), .ZN(new_n1028));
  OAI22_X1  g828(.A1(new_n729), .A2(new_n712), .B1(new_n672), .B2(new_n218), .ZN(new_n1029));
  AOI21_X1  g829(.A(new_n1029), .B1(G97), .B2(new_n665), .ZN(new_n1030));
  OAI22_X1  g830(.A1(new_n669), .A2(new_n220), .B1(new_n667), .B2(new_n315), .ZN(new_n1031));
  OAI211_X1 g831(.A(new_n341), .B(new_n280), .C1(new_n659), .C2(new_n717), .ZN(new_n1032));
  NOR2_X1   g832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g833(.A1(new_n1030), .A2(new_n887), .A3(new_n924), .A4(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g834(.A(new_n1034), .B(KEYINPUT118), .ZN(new_n1035));
  OR2_X1    g835(.A1(new_n1035), .A2(KEYINPUT58), .ZN(new_n1036));
  NAND2_X1  g836(.A1(new_n678), .A2(G125), .ZN(new_n1037));
  OAI21_X1  g837(.A(new_n1037), .B1(new_n716), .B2(new_n721), .ZN(new_n1038));
  AOI22_X1  g838(.A1(new_n670), .A2(G128), .B1(new_n725), .B2(G137), .ZN(new_n1039));
  OAI21_X1  g839(.A(new_n1039), .B1(new_n656), .B2(new_n976), .ZN(new_n1040));
  AOI211_X1 g840(.A(new_n1038), .B(new_n1040), .C1(G150), .C2(new_n677), .ZN(new_n1041));
  INV_X1    g841(.A(new_n1041), .ZN(new_n1042));
  OR2_X1    g842(.A1(new_n1042), .A2(KEYINPUT59), .ZN(new_n1043));
  NAND2_X1  g843(.A1(new_n1042), .A2(KEYINPUT59), .ZN(new_n1044));
  NAND2_X1  g844(.A1(new_n673), .A2(G159), .ZN(new_n1045));
  AOI211_X1 g845(.A(G33), .B(G41), .C1(new_n660), .C2(G124), .ZN(new_n1046));
  NAND4_X1  g846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  OAI221_X1 g847(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n450), .C2(new_n270), .ZN(new_n1048));
  NAND2_X1  g848(.A1(new_n1035), .A2(KEYINPUT58), .ZN(new_n1049));
  NAND4_X1  g849(.A1(new_n1036), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g850(.A(new_n1028), .B1(new_n1050), .B2(new_n651), .ZN(new_n1051));
  NAND2_X1  g851(.A1(new_n1027), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g852(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g853(.A(G330), .B1(new_n790), .B2(new_n782), .ZN(new_n1054));
  INV_X1    g854(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g855(.A(new_n777), .ZN(new_n1056));
  NAND2_X1  g856(.A1(new_n782), .A2(KEYINPUT102), .ZN(new_n1057));
  NAND3_X1  g857(.A1(new_n803), .A2(new_n771), .A3(new_n779), .ZN(new_n1058));
  NAND3_X1  g858(.A1(new_n1057), .A2(new_n763), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g859(.A(new_n776), .B1(new_n1059), .B2(new_n744), .ZN(new_n1060));
  OAI21_X1  g860(.A(new_n1055), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g861(.A1(new_n1061), .A2(KEYINPUT120), .ZN(new_n1062));
  INV_X1    g862(.A(KEYINPUT120), .ZN(new_n1063));
  NAND3_X1  g863(.A1(new_n778), .A2(new_n1063), .A3(new_n1055), .ZN(new_n1064));
  INV_X1    g864(.A(new_n1026), .ZN(new_n1065));
  NAND3_X1  g865(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND4_X1  g866(.A1(new_n778), .A2(new_n1063), .A3(new_n1055), .A4(new_n1026), .ZN(new_n1067));
  AND3_X1   g867(.A1(new_n1066), .A2(new_n810), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g868(.A(new_n810), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1069));
  NOR2_X1   g869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g870(.A(new_n1053), .B1(new_n1070), .B2(new_n630), .ZN(new_n1071));
  INV_X1    g871(.A(new_n1014), .ZN(new_n1072));
  NAND2_X1  g872(.A1(new_n1019), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g873(.A(KEYINPUT57), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g874(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1075));
  NAND2_X1  g875(.A1(new_n1075), .A2(new_n809), .ZN(new_n1076));
  INV_X1    g876(.A(KEYINPUT57), .ZN(new_n1077));
  AOI21_X1  g877(.A(new_n1077), .B1(new_n1019), .B2(new_n1072), .ZN(new_n1078));
  NAND3_X1  g878(.A1(new_n1066), .A2(new_n810), .A3(new_n1067), .ZN(new_n1079));
  NAND3_X1  g879(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g880(.A1(new_n1080), .A2(new_n627), .ZN(new_n1081));
  OAI21_X1  g881(.A(new_n1071), .B1(new_n1074), .B2(new_n1081), .ZN(G375));
  NAND2_X1  g882(.A1(new_n1010), .A2(new_n630), .ZN(new_n1083));
  OAI21_X1  g883(.A(new_n631), .B1(new_n707), .B2(G68), .ZN(new_n1084));
  OAI22_X1  g884(.A1(new_n712), .A2(new_n716), .B1(new_n729), .B2(new_n454), .ZN(new_n1085));
  AOI21_X1  g885(.A(new_n1085), .B1(G97), .B2(new_n688), .ZN(new_n1086));
  AOI21_X1  g886(.A(new_n270), .B1(new_n660), .B2(G303), .ZN(new_n1087));
  AOI22_X1  g887(.A1(new_n670), .A2(G283), .B1(new_n725), .B2(new_n301), .ZN(new_n1088));
  AOI22_X1  g888(.A1(new_n677), .A2(new_n922), .B1(new_n673), .B2(G77), .ZN(new_n1089));
  NAND4_X1  g889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g890(.A1(new_n678), .A2(G132), .ZN(new_n1091));
  OAI221_X1 g891(.A(new_n1091), .B1(new_n728), .B2(new_n669), .C1(new_n716), .C2(new_n976), .ZN(new_n1092));
  NOR2_X1   g892(.A1(new_n1092), .A2(KEYINPUT121), .ZN(new_n1093));
  NAND2_X1  g893(.A1(new_n1092), .A2(KEYINPUT121), .ZN(new_n1094));
  OAI21_X1  g894(.A(new_n270), .B1(new_n667), .B2(new_n727), .ZN(new_n1095));
  AOI21_X1  g895(.A(new_n1095), .B1(G128), .B2(new_n660), .ZN(new_n1096));
  OAI22_X1  g896(.A1(new_n218), .A2(new_n672), .B1(new_n656), .B2(new_n350), .ZN(new_n1097));
  AOI21_X1  g897(.A(new_n1097), .B1(G50), .B2(new_n677), .ZN(new_n1098));
  NAND3_X1  g898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g899(.A(new_n1090), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g900(.A(new_n1084), .B1(new_n1100), .B2(new_n651), .ZN(new_n1101));
  OAI21_X1  g901(.A(new_n1101), .B1(new_n803), .B2(new_n636), .ZN(new_n1102));
  NAND2_X1  g902(.A1(new_n1083), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g904(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1105));
  INV_X1    g905(.A(new_n876), .ZN(new_n1106));
  NAND2_X1  g906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g907(.A(new_n1104), .B1(new_n1016), .B2(new_n1107), .ZN(G381));
  NAND3_X1  g908(.A1(new_n910), .A2(new_n694), .A3(new_n949), .ZN(new_n1109));
  NOR3_X1   g909(.A1(G390), .A2(G384), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g910(.A1(new_n906), .A2(new_n1110), .ZN(new_n1111));
  OR4_X1    g911(.A1(G378), .A2(new_n1111), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g912(.A(G213), .ZN(new_n1113));
  NOR2_X1   g913(.A1(new_n1113), .A2(G343), .ZN(new_n1114));
  NAND2_X1  g914(.A1(new_n1020), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g915(.A(G407), .B(G213), .C1(G375), .C2(new_n1115), .ZN(G409));
  NAND2_X1  g916(.A1(G393), .A2(G396), .ZN(new_n1117));
  NAND2_X1  g917(.A1(new_n1117), .A2(new_n1109), .ZN(new_n1118));
  NAND2_X1  g918(.A1(new_n1118), .A2(KEYINPUT111), .ZN(new_n1119));
  NAND3_X1  g919(.A1(new_n1119), .A2(new_n954), .A3(new_n974), .ZN(new_n1120));
  NAND2_X1  g920(.A1(G390), .A2(new_n1118), .ZN(new_n1121));
  NAND3_X1  g921(.A1(new_n905), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  NAND3_X1  g923(.A1(new_n1123), .A2(new_n878), .A3(new_n904), .ZN(new_n1124));
  NAND2_X1  g924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g925(.A(KEYINPUT61), .ZN(new_n1126));
  OAI211_X1 g926(.A(G378), .B(new_n1071), .C1(new_n1074), .C2(new_n1081), .ZN(new_n1127));
  NAND4_X1  g927(.A1(new_n1076), .A2(new_n1106), .A3(new_n1079), .A4(new_n1073), .ZN(new_n1128));
  NAND3_X1  g928(.A1(new_n1076), .A2(new_n630), .A3(new_n1079), .ZN(new_n1129));
  NAND3_X1  g929(.A1(new_n1128), .A2(new_n1129), .A3(new_n1052), .ZN(new_n1130));
  NAND2_X1  g930(.A1(new_n1130), .A2(new_n1020), .ZN(new_n1131));
  AOI21_X1  g931(.A(new_n1114), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g932(.A1(new_n1114), .A2(G2897), .ZN(new_n1133));
  INV_X1    g933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g934(.A1(new_n1011), .A2(new_n1015), .A3(KEYINPUT60), .ZN(new_n1135));
  NAND2_X1  g935(.A1(new_n1135), .A2(new_n1105), .ZN(new_n1136));
  INV_X1    g936(.A(KEYINPUT60), .ZN(new_n1137));
  OAI21_X1  g937(.A(new_n627), .B1(new_n1105), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g940(.A1(new_n1140), .A2(G384), .A3(new_n1104), .ZN(new_n1141));
  AOI21_X1  g941(.A(new_n1138), .B1(new_n1135), .B2(new_n1105), .ZN(new_n1142));
  OAI21_X1  g942(.A(new_n734), .B1(new_n1142), .B2(new_n1103), .ZN(new_n1143));
  NAND2_X1  g943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g944(.A(new_n1134), .B1(new_n1144), .B2(KEYINPUT122), .ZN(new_n1145));
  NAND2_X1  g945(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1146));
  NAND2_X1  g946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g947(.A(new_n1147), .B1(new_n1146), .B2(new_n1133), .ZN(new_n1148));
  INV_X1    g948(.A(new_n1144), .ZN(new_n1149));
  NAND2_X1  g949(.A1(new_n1132), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g950(.A(new_n1126), .B1(new_n1132), .B2(new_n1148), .C1(new_n1150), .C2(KEYINPUT62), .ZN(new_n1151));
  AND2_X1   g951(.A1(new_n1150), .A2(KEYINPUT62), .ZN(new_n1152));
  OAI21_X1  g952(.A(new_n1125), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g953(.A1(new_n1122), .A2(new_n1126), .A3(new_n1124), .ZN(new_n1154));
  NAND2_X1  g954(.A1(new_n1154), .A2(KEYINPUT123), .ZN(new_n1155));
  INV_X1    g955(.A(KEYINPUT123), .ZN(new_n1156));
  NAND4_X1  g956(.A1(new_n1122), .A2(new_n1156), .A3(new_n1126), .A4(new_n1124), .ZN(new_n1157));
  NAND2_X1  g957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g958(.A(new_n1158), .B1(new_n1132), .B2(new_n1148), .ZN(new_n1159));
  AOI21_X1  g959(.A(KEYINPUT63), .B1(new_n1132), .B2(new_n1149), .ZN(new_n1160));
  NOR2_X1   g960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g961(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1162));
  INV_X1    g962(.A(new_n1114), .ZN(new_n1163));
  AND2_X1   g963(.A1(new_n1149), .A2(KEYINPUT63), .ZN(new_n1164));
  NAND3_X1  g964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g965(.A1(new_n1165), .A2(KEYINPUT124), .ZN(new_n1166));
  INV_X1    g966(.A(KEYINPUT124), .ZN(new_n1167));
  NAND3_X1  g967(.A1(new_n1132), .A2(new_n1167), .A3(new_n1164), .ZN(new_n1168));
  NAND2_X1  g968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g969(.A(KEYINPUT125), .ZN(new_n1170));
  AND3_X1   g970(.A1(new_n1161), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g971(.A(new_n1170), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1172));
  OAI21_X1  g972(.A(new_n1153), .B1(new_n1171), .B2(new_n1172), .ZN(G405));
  AND2_X1   g973(.A1(G375), .A2(new_n1020), .ZN(new_n1174));
  INV_X1    g974(.A(new_n1127), .ZN(new_n1175));
  NOR2_X1   g975(.A1(new_n1144), .A2(KEYINPUT126), .ZN(new_n1176));
  OR3_X1    g976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g977(.A(new_n1176), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1178));
  NAND2_X1  g978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g979(.A(new_n1179), .B(new_n1125), .ZN(G402));
endmodule


