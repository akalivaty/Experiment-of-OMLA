//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT80), .B1(new_n187), .B2(G125), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G140), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n191), .A2(new_n194), .B1(G125), .B2(new_n187), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(new_n189), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(new_n190), .C1(new_n195), .C2(new_n189), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT81), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT71), .B(G119), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G128), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT79), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n209), .B(new_n210), .C1(KEYINPUT23), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G110), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n196), .A2(new_n214), .A3(G146), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n200), .A2(new_n206), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n212), .A2(G110), .B1(new_n204), .B2(new_n205), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n193), .A2(G140), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n188), .A2(new_n218), .A3(new_n198), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n197), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n222), .B(new_n224), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n220), .A3(new_n225), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n232));
  OR3_X1    g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(G234), .B2(new_n228), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n232), .B1(new_n230), .B2(new_n231), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT83), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT83), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n239), .A3(new_n235), .A4(new_n236), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n227), .A2(new_n229), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n235), .A2(G902), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n203), .A2(G116), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n201), .A2(G116), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(KEYINPUT70), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n247), .B1(new_n203), .B2(G116), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n198), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n260), .A3(G128), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT68), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G143), .B(G146), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .A4(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n198), .A2(G143), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n273), .A2(new_n265), .A3(new_n267), .ZN(new_n274));
  AOI21_X1  g088(.A(G128), .B1(new_n258), .B2(new_n260), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT69), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n275), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n262), .A2(new_n273), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n272), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G134), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G137), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(KEYINPUT11), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n284), .B2(G137), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n287), .B(new_n289), .C1(G134), .C2(new_n282), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n290), .A2(G131), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n281), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT73), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n290), .B(G131), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT0), .A4(G128), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT64), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n269), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT0), .B(G128), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n269), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n299), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n294), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n281), .A2(new_n306), .A3(new_n286), .A4(new_n291), .ZN(new_n307));
  AND4_X1   g121(.A1(new_n257), .A2(new_n293), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n305), .A2(new_n307), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(KEYINPUT74), .A3(KEYINPUT30), .A4(new_n293), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n305), .A4(new_n307), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n299), .A2(new_n302), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n299), .A2(KEYINPUT65), .A3(new_n302), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n294), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n317), .A2(new_n294), .A3(new_n321), .A4(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n292), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n257), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n308), .B1(new_n314), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT26), .B(G101), .Z(new_n327));
  NOR2_X1   g141(.A1(G237), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G210), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT75), .B(KEYINPUT27), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n245), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  INV_X1    g148(.A(new_n308), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n323), .A2(new_n256), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n305), .A2(new_n257), .A3(new_n292), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n334), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n332), .B(KEYINPUT76), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n337), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT77), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n311), .B(KEYINPUT74), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n323), .A2(new_n324), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n256), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n335), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n332), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n308), .B1(new_n256), .B2(new_n323), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n339), .B(new_n341), .C1(new_n352), .C2(new_n334), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n245), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n309), .A2(new_n293), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n256), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n334), .B1(new_n356), .B2(new_n335), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(new_n340), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n349), .A2(new_n245), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n344), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n361), .A2(KEYINPUT78), .A3(G472), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT78), .B1(new_n361), .B2(G472), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n335), .B(new_n332), .C1(new_n345), .C2(new_n347), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT31), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n326), .A2(new_n367), .A3(new_n332), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n342), .B1(new_n337), .B2(new_n340), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT32), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n244), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  XOR2_X1   g190(.A(G110), .B(G122), .Z(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT86), .B(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(G101), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(G101), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n379), .A2(new_n382), .A3(new_n389), .A4(new_n383), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT85), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n393), .A3(KEYINPUT4), .A4(new_n390), .ZN(new_n394));
  AOI221_X4 g208(.A(new_n387), .B1(new_n251), .B2(new_n255), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n383), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n378), .A2(G107), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n390), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n253), .A2(new_n252), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G116), .ZN(new_n403));
  NOR2_X1   g217(.A1(KEYINPUT71), .A2(G119), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT71), .A2(G119), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n407), .A2(new_n408), .A3(new_n247), .ZN(new_n409));
  OAI21_X1  g223(.A(G113), .B1(new_n246), .B2(KEYINPUT5), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT87), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G113), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n407), .B2(new_n408), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(new_n414), .C1(new_n408), .C2(new_n249), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n402), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n377), .B1(new_n395), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n392), .A2(new_n394), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n256), .A3(new_n386), .ZN(new_n420));
  INV_X1    g234(.A(new_n377), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n422), .A3(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT88), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n417), .A2(new_n422), .A3(new_n425), .A4(KEYINPUT6), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT89), .B1(new_n417), .B2(KEYINPUT6), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n421), .B1(new_n418), .B2(new_n420), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n281), .A2(G125), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n315), .A2(G125), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT90), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n315), .A2(new_n437), .A3(G125), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G953), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n427), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n434), .A2(new_n438), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n445), .A2(new_n436), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n439), .A2(new_n448), .B1(new_n446), .B2(new_n441), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n377), .B(KEYINPUT8), .Z(new_n452));
  NAND2_X1  g266(.A1(new_n411), .A2(new_n415), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n400), .B1(new_n453), .B2(new_n401), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n409), .A2(new_n410), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n402), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n452), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n450), .A2(new_n451), .A3(new_n422), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n228), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n443), .A2(new_n444), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n444), .B1(new_n443), .B2(new_n460), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n376), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n200), .A2(new_n215), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n328), .A2(G143), .A3(G214), .ZN(new_n465));
  AOI21_X1  g279(.A(G143), .B1(new_n328), .B2(G214), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n468));
  INV_X1    g282(.A(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n223), .A3(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n259), .ZN(new_n471));
  INV_X1    g285(.A(G131), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n328), .A2(G143), .A3(G214), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n467), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(new_n473), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT17), .A3(G131), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n464), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n378), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n478), .B(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n219), .B1(new_n195), .B2(new_n198), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n467), .A2(new_n474), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT19), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n188), .A2(new_n218), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n195), .B2(new_n489), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n197), .B(new_n488), .C1(G146), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n486), .ZN(new_n493));
  INV_X1    g307(.A(new_n482), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(KEYINPUT92), .A3(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n487), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G475), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n228), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n499), .A2(new_n503), .A3(new_n500), .A4(new_n228), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n482), .B1(new_n480), .B2(new_n486), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT94), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n507), .B(new_n228), .C1(new_n509), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G475), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n207), .B2(G143), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n259), .A2(KEYINPUT95), .A3(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n259), .A2(G128), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n517), .A2(G134), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(G116), .B(G122), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(G107), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n524));
  INV_X1    g338(.A(new_n518), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(KEYINPUT13), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT13), .B1(new_n514), .B2(new_n515), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT96), .B1(new_n528), .B2(new_n518), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AOI211_X1 g344(.A(new_n519), .B(new_n521), .C1(new_n530), .C2(G134), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n520), .A2(new_n381), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n403), .A2(KEYINPUT14), .A3(G122), .ZN(new_n533));
  INV_X1    g347(.A(new_n520), .ZN(new_n534));
  OAI211_X1 g348(.A(G107), .B(new_n533), .C1(new_n534), .C2(KEYINPUT14), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n284), .B1(new_n516), .B2(new_n525), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n532), .B(new_n535), .C1(new_n519), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT9), .B(G234), .Z(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(G217), .A3(new_n223), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n531), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n540), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n521), .B1(new_n530), .B2(G134), .ZN(new_n543));
  INV_X1    g357(.A(new_n519), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n545), .B2(new_n537), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n228), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G478), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(KEYINPUT15), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n547), .A2(new_n549), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n512), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G469), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n263), .A2(new_n271), .B1(KEYINPUT1), .B2(new_n273), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n399), .B1(new_n555), .B2(new_n277), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n556), .A2(KEYINPUT10), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n419), .B(new_n386), .C1(new_n304), .C2(new_n303), .ZN(new_n558));
  INV_X1    g372(.A(new_n294), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n400), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n281), .A2(new_n400), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n294), .B1(new_n563), .B2(new_n556), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT12), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n294), .C1(new_n563), .C2(new_n556), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n223), .A2(G227), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n562), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n294), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n575), .B2(new_n561), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n554), .B(new_n228), .C1(new_n573), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n554), .A2(new_n228), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n572), .B1(new_n562), .B2(new_n568), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n561), .A3(new_n571), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(G469), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G221), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n539), .B2(new_n228), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT84), .Z(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n223), .A2(G952), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(G234), .B2(G237), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT21), .B(G898), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n228), .B(new_n223), .C1(G234), .C2(G237), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR4_X1   g407(.A1(new_n463), .A2(new_n553), .A3(new_n587), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n375), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  NAND2_X1  g410(.A1(new_n370), .A2(new_n228), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n597), .A2(G472), .B1(new_n371), .B2(new_n370), .ZN(new_n598));
  INV_X1    g412(.A(new_n587), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT99), .B(G478), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n547), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n545), .B2(new_n537), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  OAI22_X1  g419(.A1(new_n541), .A2(new_n546), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n540), .B1(new_n531), .B2(new_n538), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT97), .B1(new_n531), .B2(new_n538), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n545), .A2(new_n537), .A3(new_n542), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(KEYINPUT33), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n606), .A2(G478), .A3(new_n228), .A4(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n602), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n505), .A2(new_n511), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n463), .A2(new_n244), .A3(new_n593), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n600), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G104), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n552), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n512), .A2(new_n623), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n463), .A2(new_n244), .A3(new_n624), .A4(new_n593), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n600), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT35), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT101), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT102), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n221), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n242), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n238), .A2(new_n240), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n598), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(new_n594), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NAND2_X1  g454(.A1(new_n361), .A2(G472), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT78), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n361), .A2(KEYINPUT78), .A3(G472), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n374), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n634), .A2(new_n599), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n589), .B1(new_n592), .B2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n463), .A2(new_n624), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XNOR2_X1  g466(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n649), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n599), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n461), .A2(new_n462), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n657), .A2(new_n634), .A3(new_n659), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n308), .B(new_n349), .C1(new_n314), .C2(new_n325), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n369), .B1(new_n661), .B2(new_n367), .ZN(new_n662));
  INV_X1    g476(.A(new_n368), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n371), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT32), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n370), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n341), .B1(new_n356), .B2(new_n335), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n228), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G472), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n552), .B1(new_n505), .B2(new_n511), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n655), .B2(KEYINPUT40), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n660), .A2(new_n376), .A3(new_n671), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(new_n649), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n615), .A2(new_n616), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n463), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n645), .A2(new_n647), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(new_n228), .B1(new_n573), .B2(new_n576), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  INV_X1    g497(.A(new_n585), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n577), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n645), .A2(new_n618), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NOR2_X1   g503(.A1(new_n463), .A2(new_n685), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n645), .A2(new_n625), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  INV_X1    g506(.A(new_n634), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n553), .A3(new_n593), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n645), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NOR3_X1   g510(.A1(new_n463), .A2(new_n244), .A3(new_n593), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n339), .B1(new_n352), .B2(new_n334), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n365), .A2(KEYINPUT31), .B1(new_n698), .B2(new_n342), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n699), .B2(new_n368), .ZN(new_n700));
  INV_X1    g514(.A(G472), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT106), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n597), .A2(new_n703), .A3(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n673), .A2(new_n685), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n342), .B1(new_n357), .B2(new_n340), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n366), .A2(new_n368), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n371), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n708), .B2(new_n371), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n697), .A2(new_n705), .A3(new_n706), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR3_X1   g529(.A1(new_n463), .A2(new_n678), .A3(new_n685), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n705), .A2(new_n716), .A3(new_n713), .A4(new_n634), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  INV_X1    g532(.A(new_n244), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n658), .A2(new_n376), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n577), .A2(new_n579), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT107), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n575), .A2(new_n723), .A3(new_n561), .A4(new_n571), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n721), .B1(G469), .B2(new_n725), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n720), .A2(new_n585), .A3(new_n678), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n645), .A2(new_n719), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n645), .A2(new_n727), .A3(KEYINPUT42), .A4(new_n719), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  NOR2_X1   g547(.A1(new_n624), .A2(new_n649), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n720), .A2(new_n585), .A3(new_n726), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n645), .A2(new_n719), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  OR2_X1    g551(.A1(new_n611), .A2(new_n612), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n611), .A2(new_n612), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n738), .A2(new_n739), .B1(new_n547), .B2(new_n601), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n616), .A2(KEYINPUT112), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n505), .A2(new_n742), .A3(new_n511), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT43), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT43), .B1(new_n512), .B2(new_n615), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI211_X1 g562(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n512), .C2(new_n615), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n598), .A2(new_n693), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT44), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n720), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT113), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n725), .B2(KEYINPUT45), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI211_X1 g572(.A(KEYINPUT109), .B(new_n758), .C1(new_n722), .C2(new_n724), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(KEYINPUT45), .A2(G469), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n582), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n582), .A2(KEYINPUT108), .A3(new_n761), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n579), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n577), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n578), .B1(new_n760), .B2(new_n766), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(KEYINPUT46), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n772), .B2(KEYINPUT46), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(new_n684), .A3(new_n654), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT44), .B1(new_n750), .B2(new_n751), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n752), .A2(new_n780), .A3(new_n753), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n755), .A2(new_n777), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT114), .B(G137), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G39));
  NOR3_X1   g598(.A1(new_n719), .A2(new_n720), .A3(new_n678), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n364), .A2(new_n785), .A3(new_n374), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT115), .Z(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n776), .A2(new_n788), .A3(new_n684), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n788), .B1(new_n776), .B2(new_n684), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n683), .A2(new_n577), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n744), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n376), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n586), .B1(new_n795), .B2(KEYINPUT49), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n671), .A2(new_n244), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n659), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT116), .Z(new_n803));
  INV_X1    g617(.A(new_n750), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n753), .A2(new_n684), .A3(new_n589), .A4(new_n796), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n375), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n588), .B1(new_n809), .B2(KEYINPUT48), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n805), .A2(new_n244), .A3(new_n671), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n616), .A3(new_n615), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n750), .A2(new_n719), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n705), .A2(new_n713), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(new_n814), .A3(new_n589), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n690), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT48), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n807), .A2(KEYINPUT121), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n810), .A2(new_n812), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n815), .A2(new_n753), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n789), .A2(new_n790), .B1(new_n586), .B2(new_n795), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n811), .A2(new_n512), .A3(new_n740), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n806), .A2(new_n634), .A3(new_n814), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n826), .B(new_n828), .C1(new_n821), .C2(new_n822), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n813), .A2(new_n814), .A3(new_n589), .A4(new_n686), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n659), .A2(new_n798), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n830), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n824), .A2(new_n829), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n821), .A2(new_n822), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n825), .A3(new_n827), .ZN(new_n838));
  INV_X1    g652(.A(new_n835), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n838), .A2(new_n839), .B1(new_n823), .B2(KEYINPUT51), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n819), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n651), .A2(new_n680), .A3(new_n717), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n672), .B(new_n376), .C1(new_n461), .C2(new_n462), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n649), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n634), .A2(new_n726), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n671), .A2(new_n845), .A3(new_n846), .A4(new_n684), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT118), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n842), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n634), .A2(new_n705), .A3(new_n713), .A4(new_n716), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n646), .B1(new_n364), .B2(new_n374), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n851), .B2(new_n650), .ZN(new_n852));
  INV_X1    g666(.A(new_n725), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n577), .B(new_n579), .C1(new_n853), .C2(new_n554), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n240), .A3(new_n238), .A4(new_n633), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n374), .B2(new_n670), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT118), .A3(new_n684), .A4(new_n845), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n847), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n680), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n849), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n687), .A2(new_n695), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n697), .A2(new_n705), .A3(new_n706), .A4(new_n713), .ZN(new_n864));
  INV_X1    g678(.A(new_n690), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n364), .B2(new_n374), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n864), .B1(new_n866), .B2(new_n625), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n687), .A2(new_n695), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n691), .A2(new_n714), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT117), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n727), .A2(new_n634), .A3(new_n713), .A4(new_n705), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n736), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n553), .A2(new_n649), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n851), .A2(new_n753), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n732), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n595), .A2(new_n638), .A3(new_n619), .A4(new_n626), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n862), .A2(new_n873), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT53), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n869), .B2(new_n872), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n878), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n849), .B2(new_n861), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n651), .A2(new_n680), .A3(new_n717), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n860), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT119), .B1(new_n889), .B2(new_n842), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n885), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n882), .B(KEYINPUT54), .C1(new_n884), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n881), .A2(new_n885), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n732), .A2(new_n875), .A3(KEYINPUT53), .A4(new_n877), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n879), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n870), .A2(new_n871), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n895), .B(new_n896), .C1(new_n887), .C2(new_n890), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n841), .A2(new_n892), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(G952), .A2(G953), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n803), .B1(new_n900), .B2(new_n901), .ZN(G75));
  AOI22_X1  g716(.A1(new_n424), .A2(new_n426), .B1(new_n428), .B2(new_n432), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(new_n442), .Z(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  INV_X1    g719(.A(G210), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n906), .B(new_n228), .C1(new_n893), .C2(new_n897), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n907), .B2(KEYINPUT56), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  INV_X1    g723(.A(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n893), .A2(new_n897), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G902), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n909), .B(new_n910), .C1(new_n912), .C2(new_n906), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n223), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n908), .A2(new_n913), .A3(new_n915), .ZN(G51));
  XNOR2_X1  g730(.A(new_n578), .B(KEYINPUT57), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n893), .A2(new_n898), .A3(new_n897), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n898), .B1(new_n893), .B2(new_n897), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n573), .A2(new_n576), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n912), .A2(new_n767), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n922), .B2(new_n923), .ZN(G54));
  NAND2_X1  g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n911), .A2(G902), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n499), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n915), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n927), .A2(new_n932), .A3(new_n928), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n931), .B2(new_n933), .ZN(G60));
  AND2_X1   g748(.A1(new_n606), .A2(new_n610), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n935), .B(new_n937), .C1(new_n918), .C2(new_n919), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n915), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n892), .A2(new_n899), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n940), .B2(new_n937), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(G63));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n893), .B2(new_n897), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n632), .B(KEYINPUT123), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n915), .B1(new_n946), .B2(new_n241), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n241), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n893), .A2(new_n897), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n945), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT61), .A3(new_n915), .A4(new_n948), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(G66));
  OAI21_X1  g770(.A(G953), .B1(new_n591), .B2(new_n440), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n883), .B2(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n903), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(G898), .B2(new_n223), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  NAND2_X1  g775(.A1(new_n314), .A2(new_n346), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT124), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(new_n491), .ZN(new_n964));
  OAI21_X1  g778(.A(G900), .B1(new_n964), .B2(G227), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n223), .B(new_n965), .C1(G227), .C2(new_n964), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  INV_X1    g781(.A(new_n675), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n843), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n675), .A2(new_n888), .A3(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  INV_X1    g786(.A(new_n655), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n624), .A2(new_n617), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n375), .A2(new_n973), .A3(new_n753), .A4(new_n974), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n782), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n782), .B2(new_n975), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n971), .B(new_n792), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n964), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n752), .A2(new_n780), .A3(new_n753), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n780), .B1(new_n752), .B2(new_n753), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n778), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n244), .B(new_n844), .C1(new_n364), .C2(new_n374), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n777), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n888), .A2(new_n736), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n791), .B2(new_n787), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n985), .A2(new_n987), .A3(new_n732), .A4(new_n964), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n966), .B1(new_n980), .B2(new_n988), .ZN(G72));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  INV_X1    g805(.A(new_n883), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n978), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n348), .A3(new_n332), .ZN(new_n994));
  INV_X1    g808(.A(new_n991), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n350), .B2(new_n365), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n882), .B(new_n996), .C1(new_n884), .C2(new_n891), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n985), .A2(new_n987), .A3(new_n883), .A4(new_n732), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n332), .B1(new_n1000), .B2(new_n991), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n326), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n999), .B1(new_n1002), .B2(new_n915), .ZN(new_n1003));
  AOI211_X1 g817(.A(KEYINPUT126), .B(new_n914), .C1(new_n1001), .C2(new_n326), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n998), .A2(new_n1003), .A3(new_n1004), .ZN(G57));
endmodule


