//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT77), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n206), .C1(KEYINPUT22), .C2(new_n209), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G226gat), .ZN(new_n217));
  INV_X1    g016(.A(G233gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT28), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT68), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n221), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n220), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT69), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT26), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n237), .A2(new_n233), .A3(new_n234), .A4(KEYINPUT69), .ZN(new_n238));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n223), .B1(new_n245), .B2(KEYINPUT27), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n220), .A2(new_n231), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n240), .B(new_n241), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT65), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n231), .ZN(new_n255));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n251), .A2(new_n254), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G169gat), .B2(G176gat), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n258), .A2(new_n260), .A3(new_n239), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT25), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT25), .A4(new_n239), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT67), .B(G183gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n252), .B1(new_n264), .B2(new_n231), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n263), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n232), .A2(new_n248), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n219), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n219), .ZN(new_n274));
  INV_X1    g073(.A(new_n254), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n255), .B(new_n256), .C1(new_n252), .C2(new_n253), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n261), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n242), .A2(new_n244), .A3(new_n231), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(new_n250), .A3(new_n266), .A4(new_n268), .ZN(new_n281));
  INV_X1    g080(.A(new_n263), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n235), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n285), .A2(new_n238), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n225), .B1(new_n242), .B2(new_n244), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n220), .B(new_n231), .C1(new_n287), .C2(new_n223), .ZN(new_n288));
  AOI21_X1  g087(.A(G190gat), .B1(new_n224), .B2(new_n229), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n286), .B(new_n288), .C1(new_n220), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n274), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT76), .B1(new_n273), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n284), .B2(new_n290), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n219), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n216), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n271), .A2(new_n219), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n294), .B2(new_n219), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(new_n215), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n205), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n273), .A2(new_n291), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n216), .ZN(new_n302));
  INV_X1    g101(.A(new_n205), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n248), .A2(new_n232), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n277), .A2(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n272), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT76), .B1(new_n306), .B2(new_n274), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(KEYINPUT76), .B2(new_n298), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n302), .B(new_n303), .C1(new_n308), .C2(new_n216), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n300), .A2(new_n309), .A3(KEYINPUT30), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n296), .A2(new_n299), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(new_n303), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G113gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(G127gat), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G134gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n321), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n317), .B2(G120gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n319), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n331), .B(new_n332), .C1(G113gat), .C2(new_n319), .ZN(new_n333));
  OR2_X1    g132(.A1(G127gat), .A2(G134gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G127gat), .A2(G134gat), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT1), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G141gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G148gat), .ZN(new_n340));
  INV_X1    g139(.A(G148gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G155gat), .B(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT2), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(G155gat), .B2(G162gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(G155gat), .A3(G162gat), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n350), .A2(new_n351), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n340), .A2(new_n342), .B1(KEYINPUT2), .B2(new_n345), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n347), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n315), .B1(new_n338), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n322), .A2(G127gat), .A3(new_n323), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT71), .B(G127gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n327), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n363), .A2(new_n321), .B1(new_n333), .B2(new_n336), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(new_n364), .A3(KEYINPUT4), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n347), .B(new_n369), .C1(new_n356), .C2(new_n357), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n370), .A3(new_n338), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n366), .A2(KEYINPUT5), .A3(new_n367), .A4(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n359), .A3(new_n365), .A4(new_n367), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n360), .A2(new_n364), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n338), .A2(new_n358), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n367), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n378), .A3(new_n383), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n379), .A2(KEYINPUT80), .A3(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n388), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT6), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n314), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n213), .B2(new_n214), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n358), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n370), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n215), .B1(new_n402), .B2(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n403), .B(new_n399), .C1(new_n400), .C2(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(G22gat), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT82), .ZN(new_n408));
  XOR2_X1   g207(.A(G78gat), .B(G106gat), .Z(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT31), .B(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT64), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n364), .B1(new_n304), .B2(new_n305), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n284), .A2(new_n290), .A3(new_n338), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT34), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(new_n420), .A3(new_n422), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT32), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G15gat), .B(G43gat), .Z(new_n432));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n428), .B(KEYINPUT32), .C1(new_n430), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n423), .A2(new_n418), .A3(new_n424), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n427), .A2(new_n435), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n437), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n422), .ZN(new_n441));
  INV_X1    g240(.A(new_n420), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n424), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n442), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT34), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n438), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n408), .A2(new_n415), .A3(new_n407), .A4(new_n411), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n417), .A2(new_n439), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT35), .B1(new_n396), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n439), .B2(new_n448), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n440), .B2(new_n447), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n313), .A2(new_n310), .B1(new_n392), .B2(new_n394), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n417), .A2(new_n449), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n371), .A2(new_n359), .A3(new_n365), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(G225gat), .A3(G233gat), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n464), .A2(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n376), .A2(new_n367), .A3(new_n375), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(KEYINPUT39), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n384), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n393), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n310), .A2(new_n470), .A3(new_n313), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n458), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT84), .B(KEYINPUT37), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n302), .B(new_n475), .C1(new_n308), .C2(new_n216), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n301), .B2(new_n215), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n308), .B2(new_n215), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n480), .A4(new_n205), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n481), .A2(new_n392), .A3(new_n394), .A4(new_n309), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT85), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n311), .A2(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n476), .A2(new_n205), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n482), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n484), .C2(new_n485), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n474), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n396), .A2(new_n458), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT75), .B(new_n491), .C1(new_n453), .C2(new_n455), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n439), .A2(new_n448), .A3(KEYINPUT36), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n440), .A2(new_n447), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n427), .A2(new_n438), .B1(new_n435), .B2(new_n437), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT74), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n454), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT75), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n490), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n489), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n456), .B2(KEYINPUT36), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(new_n493), .A3(new_n492), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(KEYINPUT83), .A3(new_n490), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n462), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(KEYINPUT86), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  AND2_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT15), .B1(new_n508), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT87), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n515), .A2(KEYINPUT15), .A3(new_n508), .A4(new_n517), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT17), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n528), .B(new_n529), .C1(G1gat), .C2(new_n526), .ZN(new_n530));
  NOR2_X1   g329(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n534), .A4(new_n536), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n524), .B(new_n535), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT11), .B(G169gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT12), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n539), .A2(new_n552), .A3(new_n540), .A4(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT94), .B(G85gat), .Z(new_n556));
  INV_X1    g355(.A(G92gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT7), .ZN(new_n560));
  INV_X1    g359(.A(G99gat), .ZN(new_n561));
  INV_X1    g360(.A(G106gat), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT8), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n564), .B(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT95), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n525), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n568), .ZN(new_n572));
  AND2_X1   g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n572), .A2(new_n524), .B1(KEYINPUT41), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  OR2_X1    g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(KEYINPUT90), .ZN(new_n590));
  INV_X1    g389(.A(G57gat), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n591), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(G64gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT91), .B1(new_n591), .B2(G64gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n585), .B1(new_n586), .B2(new_n588), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n589), .A2(KEYINPUT90), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT20), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n532), .B1(new_n599), .B2(new_n598), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT93), .ZN(new_n607));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G183gat), .B(G211gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n605), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n584), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n570), .A2(new_n568), .B1(new_n590), .B2(new_n597), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n569), .A2(new_n598), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n590), .A4(new_n597), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT96), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  OR3_X1    g423(.A1(new_n616), .A2(new_n623), .A3(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n507), .A2(new_n555), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n395), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  INV_X1    g438(.A(new_n314), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  AND3_X1   g440(.A1(new_n636), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(KEYINPUT97), .ZN(new_n645));
  INV_X1    g444(.A(new_n636), .ZN(new_n646));
  OAI21_X1  g445(.A(G8gat), .B1(new_n646), .B2(new_n314), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n642), .B1(new_n647), .B2(KEYINPUT42), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n644), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT98), .ZN(G1325gat));
  OR3_X1    g449(.A1(new_n646), .A2(G15gat), .A3(new_n498), .ZN(new_n651));
  OAI21_X1  g450(.A(G15gat), .B1(new_n646), .B2(new_n505), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(G1326gat));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n458), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n500), .A2(new_n501), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n486), .A2(new_n483), .ZN(new_n658));
  INV_X1    g457(.A(new_n482), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n488), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n473), .A3(new_n472), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n506), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n461), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n612), .A2(new_n633), .ZN(new_n664));
  AND4_X1   g463(.A1(new_n554), .A2(new_n663), .A3(new_n584), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n516), .A3(new_n637), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT45), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n583), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n451), .A2(new_n460), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n451), .B2(new_n460), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n661), .A2(new_n505), .A3(new_n490), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n583), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI22_X1  g475(.A1(new_n507), .A2(new_n670), .B1(new_n676), .B2(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n664), .A2(new_n554), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT100), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n669), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n500), .A2(new_n489), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n461), .A2(KEYINPUT99), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n451), .A2(new_n460), .A3(new_n671), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n584), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n668), .ZN(new_n687));
  INV_X1    g486(.A(new_n678), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n680), .A2(new_n681), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n395), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n667), .A2(new_n691), .ZN(G1328gat));
  NAND3_X1  g491(.A1(new_n665), .A2(new_n512), .A3(new_n640), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT46), .Z(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n690), .B2(new_n314), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1329gat));
  NOR2_X1   g495(.A1(new_n677), .A2(new_n678), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G43gat), .B1(new_n698), .B2(new_n505), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n498), .A2(G43gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n665), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n505), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n679), .A2(new_n703), .A3(new_n689), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(KEYINPUT101), .B1(new_n665), .B2(new_n700), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n707), .A3(G43gat), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT102), .B(KEYINPUT47), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n708), .A3(new_n701), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n702), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT103), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n717), .B(new_n702), .C1(new_n709), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1330gat));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  OAI21_X1  g519(.A(G50gat), .B1(new_n698), .B2(new_n473), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n473), .A2(G50gat), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT104), .Z(new_n723));
  AND2_X1   g522(.A1(new_n665), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n720), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n720), .B(G50gat), .C1(new_n690), .C2(new_n473), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n724), .B1(KEYINPUT105), .B2(KEYINPUT48), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(G1331gat));
  NAND2_X1  g528(.A1(new_n674), .A2(new_n675), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n584), .A2(new_n613), .A3(new_n554), .A4(new_n634), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n395), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n591), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n314), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  INV_X1    g538(.A(new_n732), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n498), .B(KEYINPUT106), .ZN(new_n741));
  AOI21_X1  g540(.A(G71gat), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n703), .A2(G71gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n458), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g547(.A1(new_n676), .A2(new_n555), .A3(new_n613), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n749), .A2(KEYINPUT51), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(KEYINPUT51), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(new_n634), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n637), .A3(new_n556), .ZN(new_n753));
  NOR4_X1   g552(.A1(new_n677), .A2(new_n554), .A3(new_n612), .A4(new_n634), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n395), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n756), .B2(new_n556), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n752), .A2(new_n557), .A3(new_n640), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT109), .ZN(new_n759));
  OAI21_X1  g558(.A(G92gat), .B1(new_n755), .B2(new_n314), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(KEYINPUT108), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n759), .B(new_n762), .C1(new_n760), .C2(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n760), .B(new_n758), .C1(KEYINPUT108), .C2(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n755), .B2(new_n505), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n561), .A3(new_n456), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1338gat));
  OAI21_X1  g568(.A(G106gat), .B1(new_n755), .B2(new_n473), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n562), .A3(new_n458), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g572(.A1(new_n614), .A2(new_n555), .A3(new_n634), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n534), .B1(new_n533), .B2(new_n536), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n541), .A2(new_n543), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n549), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n553), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n634), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n622), .B1(new_n618), .B2(new_n619), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n629), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n618), .A2(new_n622), .A3(new_n619), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n624), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n782), .A2(new_n783), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n789), .B2(new_n785), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(new_n792), .B1(new_n551), .B2(new_n553), .ZN(new_n793));
  INV_X1    g592(.A(new_n632), .ZN(new_n794));
  INV_X1    g593(.A(new_n784), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n786), .A2(new_n787), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n785), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n798), .B2(KEYINPUT55), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n781), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n584), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n632), .B1(new_n791), .B2(new_n792), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n798), .A2(KEYINPUT55), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n583), .A2(new_n802), .A3(new_n780), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n613), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n776), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n458), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n498), .A2(new_n640), .A3(new_n395), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n555), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT112), .Z(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n637), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n813), .A2(new_n640), .A3(new_n450), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n317), .A3(new_n554), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1340gat));
  NOR3_X1   g615(.A1(new_n810), .A2(new_n319), .A3(new_n634), .ZN(new_n817));
  AOI21_X1  g616(.A(G120gat), .B1(new_n814), .B2(new_n633), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(G1341gat));
  OAI21_X1  g618(.A(new_n362), .B1(new_n810), .B2(new_n613), .ZN(new_n820));
  INV_X1    g619(.A(new_n362), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n821), .A3(new_n612), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT113), .Z(G1342gat));
  NAND4_X1  g623(.A1(new_n814), .A2(new_n322), .A3(new_n323), .A4(new_n584), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n810), .B2(new_n583), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G1343gat));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n703), .A2(new_n473), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n314), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n555), .A2(G141gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n640), .A2(new_n395), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n505), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n807), .B2(new_n473), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n554), .B1(KEYINPUT55), .B2(new_n798), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n843), .A2(new_n802), .B1(new_n634), .B2(new_n780), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n584), .B1(new_n844), .B2(KEYINPUT114), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n800), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n804), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n776), .B1(new_n612), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n473), .A2(new_n841), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n840), .B1(new_n842), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(new_n554), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n838), .B1(new_n339), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT117), .Z(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n854), .B(new_n857), .ZN(G1344gat));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n341), .A3(new_n633), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT118), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n505), .A2(new_n633), .A3(new_n839), .ZN(new_n862));
  INV_X1    g661(.A(new_n774), .ZN(new_n863));
  OR4_X1    g662(.A1(new_n583), .A2(new_n802), .A3(new_n780), .A4(new_n803), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n583), .B1(new_n800), .B2(new_n846), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT114), .B(new_n781), .C1(new_n793), .C2(new_n799), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n612), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n841), .B1(new_n871), .B2(new_n473), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n872), .A2(KEYINPUT120), .B1(new_n806), .B2(new_n850), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n613), .B1(new_n848), .B2(KEYINPUT119), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n867), .A2(new_n868), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n774), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n876), .B2(new_n458), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n862), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n341), .B1(new_n880), .B2(KEYINPUT121), .ZN(new_n881));
  INV_X1    g680(.A(new_n862), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n806), .A2(new_n850), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n877), .B2(new_n878), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n861), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n341), .C1(new_n852), .C2(new_n633), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n860), .B1(new_n889), .B2(new_n890), .ZN(G1345gat));
  NAND3_X1  g690(.A1(new_n836), .A2(new_n348), .A3(new_n612), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n852), .A2(new_n612), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n348), .ZN(G1346gat));
  NAND3_X1  g693(.A1(new_n836), .A2(new_n349), .A3(new_n584), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n852), .A2(new_n584), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n349), .ZN(G1347gat));
  NOR4_X1   g696(.A1(new_n807), .A2(new_n637), .A3(new_n314), .A4(new_n450), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n233), .A3(new_n554), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT122), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n637), .A2(new_n314), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n741), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT123), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n808), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n555), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(G1348gat));
  OAI21_X1  g705(.A(G176gat), .B1(new_n904), .B2(new_n634), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n898), .A2(new_n234), .A3(new_n633), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  OAI21_X1  g708(.A(new_n245), .B1(new_n904), .B2(new_n613), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n898), .A2(new_n230), .A3(new_n612), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(KEYINPUT125), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT125), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n913), .A2(KEYINPUT124), .A3(new_n914), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n912), .B2(KEYINPUT60), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n915), .A2(new_n916), .B1(new_n917), .B2(new_n919), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n904), .B2(new_n583), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT61), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n231), .A3(new_n584), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  AND4_X1   g723(.A1(new_n395), .A2(new_n806), .A3(new_n640), .A4(new_n834), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT126), .B(G197gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n554), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n505), .A2(new_n901), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n884), .B2(new_n885), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n555), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n926), .ZN(G1352gat));
  OAI21_X1  g730(.A(G204gat), .B1(new_n929), .B2(new_n634), .ZN(new_n932));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n933), .A3(new_n633), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT62), .Z(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n925), .A2(new_n207), .A3(new_n612), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n612), .B(new_n928), .C1(new_n884), .C2(new_n885), .ZN(new_n939));
  AND4_X1   g738(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n207), .B1(KEYINPUT127), .B2(new_n941), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n939), .A2(new_n942), .B1(new_n938), .B2(KEYINPUT63), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n937), .B1(new_n940), .B2(new_n943), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n929), .B2(new_n583), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n925), .A2(new_n208), .A3(new_n584), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1355gat));
endmodule


