//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1190, new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT66), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n471), .B(KEYINPUT67), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT68), .Z(new_n484));
  NOR2_X1   g059(.A1(new_n481), .A2(new_n467), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n480), .B(new_n484), .C1(G124), .C2(new_n485), .ZN(G162));
  NOR2_X1   g061(.A1(new_n467), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT69), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n467), .C1(new_n496), .C2(new_n462), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n471), .A2(G138), .A3(new_n467), .A4(new_n499), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n471), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n495), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n489), .A2(new_n494), .B1(new_n471), .B2(new_n503), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n508), .A2(KEYINPUT71), .A3(new_n501), .A4(new_n502), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n522), .B1(new_n512), .B2(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT6), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n516), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n523), .B2(new_n525), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(G88), .B1(G50), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n520), .A2(new_n521), .A3(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n516), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n529), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n516), .A2(G89), .A3(new_n526), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT77), .B(G90), .Z(new_n543));
  NAND3_X1  g118(.A1(new_n516), .A2(new_n543), .A3(new_n526), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT76), .B(G52), .Z(new_n545));
  NAND3_X1  g120(.A1(new_n545), .A2(new_n526), .A3(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n542), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n514), .A2(new_n515), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT75), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n553), .B1(new_n514), .B2(new_n515), .ZN(new_n556));
  INV_X1    g131(.A(new_n551), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n558), .A3(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n550), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  XNOR2_X1  g136(.A(KEYINPUT79), .B(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n527), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n526), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n512), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n529), .A2(new_n575), .A3(G53), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n575), .B1(new_n529), .B2(G53), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n516), .A2(new_n526), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n579), .A2(new_n512), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  NAND2_X1  g159(.A1(new_n529), .A2(G49), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n516), .A2(G74), .ZN(new_n589));
  AOI22_X1  g164(.A1(G651), .A2(new_n589), .B1(new_n527), .B2(G87), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n512), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n581), .A2(new_n594), .B1(new_n565), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n593), .A2(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n512), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n529), .A2(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n581), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND3_X1  g179(.A1(new_n516), .A2(G92), .A3(new_n526), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n552), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT81), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n614), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g190(.A(new_n614), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n583), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n583), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n471), .A2(new_n468), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2100), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n482), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n485), .A2(G123), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n653), .A2(new_n654), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n661), .B(new_n665), .Z(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT83), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(G229));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(G23), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT33), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G22), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G166), .B2(G16), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(G1971), .Z(new_n696));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n593), .A2(new_n596), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n690), .A2(new_n692), .ZN(new_n702));
  AND4_X1   g277(.A1(new_n693), .A2(new_n696), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G25), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n467), .A2(G107), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n485), .A2(G119), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n482), .A2(G131), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n708), .B1(new_n715), .B2(new_n707), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n688), .A2(G24), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n603), .B2(new_n688), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT84), .B(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n705), .A2(new_n706), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n482), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n485), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT26), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n730), .A2(new_n731), .B1(G105), .B2(new_n468), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n726), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT90), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G29), .B2(G32), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT91), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT24), .B(G34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(new_n707), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT89), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n476), .B2(new_n707), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2084), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n688), .A2(G19), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT87), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n569), .B2(new_n688), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1341), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n707), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n467), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n482), .B2(G139), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(new_n707), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G2072), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n744), .A2(new_n748), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n688), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n688), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n707), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n707), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n760), .A2(G1966), .B1(G2078), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n739), .B(new_n764), .C1(new_n737), .C2(new_n736), .ZN(new_n765));
  NAND2_X1  g340(.A1(G162), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G29), .B2(G35), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT29), .B(G2090), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT94), .B(G28), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(new_n707), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n770), .B1(new_n772), .B2(new_n774), .C1(new_n634), .C2(new_n707), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n707), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n482), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n485), .A2(G128), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT88), .B1(G104), .B2(G2105), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(KEYINPUT88), .A2(G104), .A3(G2105), .ZN(new_n783));
  OAI221_X1 g358(.A(G2104), .B1(G116), .B2(new_n467), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n779), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n688), .A2(G20), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT23), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G299), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n769), .A2(new_n776), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n762), .A2(G2078), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n688), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n688), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT96), .B(G1961), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n793), .B(new_n797), .C1(new_n767), .C2(new_n768), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n760), .A2(G1966), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  NOR2_X1   g375(.A1(G4), .A2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT86), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n613), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n765), .A2(new_n792), .A3(new_n798), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n725), .A2(new_n807), .ZN(G311));
  NAND2_X1  g383(.A1(new_n725), .A2(new_n807), .ZN(G150));
  NAND2_X1  g384(.A1(new_n527), .A2(G93), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT97), .B(G55), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n529), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n512), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G860), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n820), .A3(new_n816), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT98), .B1(new_n813), .B2(new_n815), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n814), .A2(new_n512), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n823), .A2(new_n820), .A3(new_n810), .A4(new_n812), .ZN(new_n824));
  OAI221_X1 g399(.A(new_n563), .B1(new_n564), .B2(new_n565), .C1(new_n512), .C2(new_n567), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n613), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT99), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n817), .B1(new_n830), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n819), .B1(new_n833), .B2(new_n834), .ZN(G145));
  NOR2_X1   g410(.A1(new_n733), .A2(new_n754), .ZN(new_n836));
  INV_X1    g411(.A(new_n734), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n754), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n714), .B(KEYINPUT101), .ZN(new_n839));
  INV_X1    g414(.A(new_n627), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n785), .B(new_n505), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n482), .A2(G142), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n485), .A2(G130), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n467), .A2(KEYINPUT100), .A3(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT100), .B1(new_n467), .B2(G118), .ZN(new_n846));
  OR2_X1    g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(G2104), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n842), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n841), .A2(new_n850), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n838), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n838), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n476), .B(new_n634), .ZN(new_n858));
  XOR2_X1   g433(.A(G162), .B(new_n858), .Z(new_n859));
  NAND3_X1  g434(.A1(new_n854), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n859), .B1(new_n854), .B2(new_n857), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n863), .A2(KEYINPUT40), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT40), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(G395));
  XNOR2_X1  g443(.A(new_n622), .B(new_n827), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n612), .A2(new_n583), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n607), .B(new_n611), .C1(new_n578), .C2(new_n582), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(G299), .A2(KEYINPUT102), .A3(new_n607), .A4(new_n611), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n870), .A2(new_n872), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n869), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n869), .A2(KEYINPUT103), .A3(new_n876), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n879), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n603), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n603), .B(KEYINPUT104), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n687), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G303), .B(new_n698), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G303), .B(G305), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n891), .A3(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n879), .A2(new_n885), .A3(new_n900), .A4(new_n886), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n888), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n888), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n816), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n816), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n896), .A2(new_n898), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n537), .A2(KEYINPUT105), .A3(new_n538), .A4(new_n539), .ZN(new_n909));
  INV_X1    g484(.A(new_n549), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n559), .B(new_n909), .C1(new_n910), .C2(new_n547), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT106), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n550), .A2(new_n913), .A3(new_n559), .A4(new_n909), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g490(.A1(G286), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n912), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n912), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n827), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n914), .ZN(new_n920));
  INV_X1    g495(.A(new_n916), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n821), .A2(new_n826), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n912), .A2(new_n914), .A3(new_n916), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(new_n925), .A3(new_n876), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n884), .B1(new_n919), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n908), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n917), .A2(new_n918), .A3(new_n827), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n899), .B(new_n926), .C1(new_n932), .C2(new_n884), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n933), .A3(new_n861), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n927), .A2(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n938), .B2(new_n899), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n881), .B1(new_n919), .B2(new_n925), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n908), .B1(new_n940), .B2(new_n876), .ZN(new_n941));
  AOI211_X1 g516(.A(new_n881), .B(new_n880), .C1(new_n919), .C2(new_n925), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT108), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n875), .B1(new_n932), .B2(new_n881), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  INV_X1    g520(.A(new_n880), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .A4(new_n908), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n939), .A2(new_n943), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n934), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n951));
  AND4_X1   g526(.A1(new_n907), .A2(new_n937), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n939), .A2(new_n943), .A3(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n939), .A2(new_n949), .A3(new_n929), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n952), .B1(new_n959), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g535(.A1(G303), .A2(G8), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(KEYINPUT113), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n496), .A2(new_n462), .ZN(new_n969));
  INV_X1    g544(.A(G125), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n473), .ZN(new_n972));
  OAI21_X1  g547(.A(G2105), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(G40), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(G1384), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n505), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n507), .B2(new_n509), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT110), .B(new_n978), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT111), .B(G1971), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n510), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT112), .B(G2090), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n505), .A2(new_n987), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n975), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n985), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT116), .B(new_n968), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n698), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n998), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n990), .A2(new_n975), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n994), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1007), .B(new_n1004), .C1(new_n1006), .C2(G288), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1006), .B2(G288), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n505), .A2(new_n986), .A3(new_n987), .ZN(new_n1012));
  INV_X1    g587(.A(G40), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n470), .A2(new_n474), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n501), .A2(new_n502), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT71), .B1(new_n1016), .B2(new_n508), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n505), .A2(new_n506), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n987), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n989), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n994), .B1(new_n985), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1011), .B1(new_n1022), .B2(new_n967), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n994), .B1(new_n985), .B2(new_n992), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n967), .ZN(new_n1026));
  INV_X1    g601(.A(G1966), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n975), .B1(new_n990), .B2(new_n976), .ZN(new_n1028));
  INV_X1    g603(.A(new_n977), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n507), .B2(new_n509), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1030), .B2(KEYINPUT117), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1032), .B(new_n1029), .C1(new_n507), .C2(new_n509), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1027), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1035));
  INV_X1    g610(.A(G2084), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1035), .B(new_n1036), .C1(new_n986), .C2(new_n979), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n994), .B(G286), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n995), .A2(new_n1023), .A3(new_n1026), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(KEYINPUT118), .A3(new_n1040), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1022), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n968), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n1023), .A3(KEYINPUT63), .A4(new_n1038), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(G301), .B(KEYINPUT54), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n982), .A2(new_n983), .ZN(new_n1051));
  INV_X1    g626(.A(G2078), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT126), .B1(new_n1020), .B2(G1961), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1035), .B1(new_n979), .B2(new_n986), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT126), .ZN(new_n1056));
  INV_X1    g631(.A(G1961), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n505), .A2(new_n977), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1052), .A2(KEYINPUT53), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1028), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1054), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1050), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1064), .A2(new_n1060), .B1(new_n1057), .B2(new_n1055), .ZN(new_n1065));
  AOI21_X1  g640(.A(G2078), .B1(new_n982), .B2(new_n983), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1065), .B(new_n1049), .C1(KEYINPUT53), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n1026), .A3(new_n1023), .A4(new_n995), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1034), .A2(G168), .A3(new_n1037), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(G168), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT51), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1075), .A3(G8), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1069), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n583), .B(KEYINPUT57), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n988), .A2(new_n991), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g660(.A(KEYINPUT119), .B(G1956), .C1(new_n988), .C2(new_n991), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n978), .B(new_n1088), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1081), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT50), .B(G1384), .C1(new_n507), .C2(new_n509), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1014), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1084), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT119), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1083), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1019), .A2(new_n976), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(new_n1090), .A3(new_n978), .A4(new_n1088), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1089), .A2(KEYINPUT120), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1098), .A2(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1080), .ZN(new_n1104));
  INV_X1    g679(.A(G2067), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1055), .A2(new_n804), .B1(new_n1105), .B2(new_n1003), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n614), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1093), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1103), .B2(new_n1080), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1087), .A2(new_n1091), .A3(new_n1081), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1092), .B2(new_n1109), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1092), .A2(new_n1104), .A3(KEYINPUT61), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1106), .B2(KEYINPUT60), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(new_n614), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1003), .A2(new_n1105), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT60), .B(new_n1121), .C1(new_n1020), .C2(G1348), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT124), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1106), .A2(new_n1118), .A3(KEYINPUT60), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n613), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT121), .B(G1996), .Z(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n980), .A2(new_n1127), .B1(new_n1003), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n569), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT59), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1116), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1108), .B1(new_n1115), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1079), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n995), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1053), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1138), .A2(new_n1065), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1137), .A2(G301), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT125), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT62), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1136), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n1045), .A2(new_n968), .A3(new_n1011), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1004), .B(KEYINPUT114), .Z(new_n1147));
  AND3_X1   g722(.A1(new_n1005), .A2(new_n1006), .A3(new_n687), .ZN(new_n1148));
  INV_X1    g723(.A(new_n998), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT115), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1146), .A2(new_n1153), .A3(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1048), .A2(new_n1134), .A3(new_n1145), .A4(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n785), .B(new_n1105), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n733), .A2(G1996), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1157), .B(new_n1158), .C1(new_n837), .C2(G1996), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n714), .B(new_n717), .Z(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n603), .B(G1986), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n990), .A2(new_n976), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n975), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1156), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1165), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(G1996), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT46), .Z(new_n1170));
  INV_X1    g745(.A(new_n1157), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1165), .B1(new_n1171), .B2(new_n733), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1168), .A2(G1986), .A3(G290), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT48), .Z(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1161), .B2(new_n1168), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n715), .A2(new_n717), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT127), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1159), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n785), .A2(G2067), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1165), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1174), .A2(new_n1177), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1167), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g759(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1186));
  OAI21_X1  g760(.A(new_n1186), .B1(new_n864), .B2(new_n862), .ZN(new_n1187));
  AND2_X1   g761(.A1(new_n937), .A2(new_n951), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n950), .B2(new_n1188), .ZN(G308));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n950), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n863), .A2(new_n865), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n1190), .A2(new_n1191), .A3(new_n1186), .ZN(G225));
endmodule


