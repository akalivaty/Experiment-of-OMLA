//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT71), .B(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n206), .B2(new_n207), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n215), .A2(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT25), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n217), .A2(new_n223), .A3(new_n229), .A4(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  OR3_X1    g032(.A1(new_n233), .A2(new_n213), .A3(KEYINPUT66), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n233), .B2(new_n213), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  INV_X1    g035(.A(new_n213), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT26), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n213), .A2(KEYINPUT67), .A3(new_n239), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n234), .A2(new_n235), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G183gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT27), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(KEYINPUT65), .B2(KEYINPUT28), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT27), .B(G183gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(G190gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n251), .A2(new_n253), .B1(KEYINPUT65), .B2(KEYINPUT28), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n219), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n232), .B1(new_n241), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n255), .A2(new_n241), .A3(KEYINPUT68), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n247), .B1(new_n246), .B2(new_n249), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n251), .A2(KEYINPUT65), .A3(KEYINPUT28), .A4(new_n248), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n262), .A2(new_n263), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n234), .A2(new_n235), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n240), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n261), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n232), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n258), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n259), .B1(new_n271), .B2(KEYINPUT72), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT68), .B1(new_n255), .B2(new_n241), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n264), .A2(new_n267), .A3(new_n261), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n231), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n257), .B1(new_n275), .B2(KEYINPUT29), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n212), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n258), .A2(KEYINPUT29), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n256), .A2(new_n280), .B1(new_n275), .B2(new_n258), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(new_n212), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G8gat), .B(G36gat), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT73), .ZN(new_n285));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT76), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G141gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(G148gat), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n292), .A2(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  OR2_X1    g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(KEYINPUT2), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  AND2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT74), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n304), .B(new_n307), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n291), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n302), .A2(new_n291), .A3(new_n310), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT3), .A3(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G127gat), .B(G134gat), .Z(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(KEYINPUT1), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G113gat), .B(G120gat), .Z(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n310), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n317), .A2(new_n321), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n327), .A2(KEYINPUT4), .A3(new_n302), .A4(new_n310), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(new_n323), .B2(new_n322), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n326), .A2(new_n332), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n302), .A2(new_n291), .A3(new_n310), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(new_n311), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n324), .B1(new_n338), .B2(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n328), .A2(new_n330), .A3(new_n333), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n323), .A2(new_n322), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n338), .B2(new_n322), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(new_n333), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n336), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT0), .ZN(new_n347));
  XNOR2_X1  g146(.A(G57gat), .B(G85gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n336), .B(new_n349), .C1(new_n341), .C2(new_n344), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n351), .A2(KEYINPUT78), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(KEYINPUT6), .A3(new_n350), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT6), .B1(new_n345), .B2(new_n350), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT78), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n290), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n279), .A2(KEYINPUT30), .A3(new_n283), .A4(new_n287), .ZN(new_n360));
  INV_X1    g159(.A(new_n287), .ZN(new_n361));
  INV_X1    g160(.A(new_n212), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n276), .A2(new_n277), .B1(new_n258), .B2(new_n256), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n271), .A2(KEYINPUT72), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n365), .B2(new_n282), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n202), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n355), .A3(new_n354), .ZN(new_n372));
  INV_X1    g171(.A(new_n367), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT79), .A4(new_n290), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n269), .A2(new_n322), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n275), .A2(new_n327), .ZN(new_n377));
  INV_X1    g176(.A(G227gat), .ZN(new_n378));
  INV_X1    g177(.A(G233gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n382), .B(KEYINPUT34), .Z(new_n383));
  XNOR2_X1  g182(.A(G15gat), .B(G43gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n275), .A2(new_n327), .ZN(new_n387));
  AOI211_X1 g186(.A(new_n322), .B(new_n231), .C1(new_n273), .C2(new_n274), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n381), .B1(new_n376), .B2(new_n377), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT70), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT70), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n395), .A3(KEYINPUT32), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n389), .B(KEYINPUT32), .C1(new_n390), .C2(new_n386), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n383), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n383), .B1(new_n397), .B2(new_n398), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G228gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n379), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n270), .B1(new_n323), .B2(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n212), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n206), .A2(new_n207), .ZN(new_n412));
  INV_X1    g211(.A(new_n208), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n414), .B2(new_n209), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n415), .B2(KEYINPUT80), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n270), .B1(new_n210), .B2(new_n211), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n323), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n410), .B1(new_n420), .B2(KEYINPUT81), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT3), .B1(new_n417), .B2(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n415), .A2(KEYINPUT80), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n422), .A2(new_n423), .B1(new_n302), .B2(new_n310), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n407), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n338), .B1(KEYINPUT3), .B2(new_n415), .ZN(new_n428));
  INV_X1    g227(.A(new_n407), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n408), .B2(new_n212), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n428), .A2(KEYINPUT82), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT82), .B1(new_n428), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(G22gat), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n427), .A2(G22gat), .A3(new_n433), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n409), .B1(new_n424), .B2(new_n425), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n420), .A2(KEYINPUT81), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n429), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n433), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n438), .A3(new_n442), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT83), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n405), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n421), .A2(new_n426), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n433), .B1(new_n448), .B2(new_n429), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n404), .B1(new_n449), .B2(new_n438), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(G22gat), .C1(new_n427), .C2(new_n433), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n447), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n401), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT35), .B1(new_n375), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n401), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(KEYINPUT83), .B2(new_n444), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n449), .A2(new_n436), .A3(new_n438), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n404), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n447), .A2(new_n450), .A3(new_n452), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n373), .A2(new_n290), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n369), .A2(new_n355), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(KEYINPUT35), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n399), .B2(new_n400), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n397), .A2(new_n398), .ZN(new_n468));
  INV_X1    g267(.A(new_n383), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n383), .A2(new_n397), .A3(new_n398), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT36), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n446), .A2(new_n453), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n375), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n212), .B1(new_n363), .B2(new_n364), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT37), .B1(new_n281), .B2(new_n362), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n361), .A2(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n366), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n288), .A2(new_n369), .A3(new_n355), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT86), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n362), .B1(new_n272), .B2(new_n278), .ZN(new_n484));
  INV_X1    g283(.A(new_n478), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n279), .A2(new_n283), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n486), .B(new_n361), .C1(KEYINPUT37), .C2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n288), .A2(new_n369), .A3(new_n355), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n487), .A2(KEYINPUT37), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n361), .B1(new_n487), .B2(KEYINPUT37), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n483), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n459), .A2(new_n460), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n343), .A2(new_n333), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT39), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n333), .B1(new_n326), .B2(new_n332), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(new_n350), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(KEYINPUT40), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT40), .B1(new_n501), .B2(new_n503), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n345), .B2(new_n350), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n462), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n495), .A2(new_n496), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n455), .A2(new_n465), .B1(new_n475), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT14), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT15), .B1(new_n518), .B2(G50gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n518), .B2(G50gat), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n517), .B(new_n520), .C1(G29gat), .C2(G36gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n518), .A2(G50gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT88), .B(G50gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n524), .B2(new_n518), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n517), .A2(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n528), .B2(new_n517), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n520), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT90), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n527), .A2(KEYINPUT17), .A3(new_n531), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT16), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(G1gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(G1gat), .B2(new_n542), .ZN(new_n545));
  INV_X1    g344(.A(G8gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n538), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n549), .A4(new_n551), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n532), .B(new_n550), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n549), .B(KEYINPUT13), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G197gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT12), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n552), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n555), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n511), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT93), .ZN(new_n574));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(KEYINPUT95), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(KEYINPUT95), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(G85gat), .B2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT96), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT94), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n583), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT97), .B1(new_n589), .B2(new_n591), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n538), .B(new_n541), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n591), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n532), .A3(new_n592), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n600), .A2(KEYINPUT98), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n577), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n576), .A3(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n615));
  XNOR2_X1  g414(.A(G57gat), .B(G64gat), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G71gat), .B(G78gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n589), .A2(new_n620), .A3(new_n591), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n589), .B2(new_n591), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n614), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n620), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n625), .A4(new_n592), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n613), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n622), .A2(new_n612), .A3(new_n623), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630));
  XOR2_X1   g429(.A(G120gat), .B(G148gat), .Z(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(KEYINPUT10), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n593), .A2(new_n594), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n614), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n596), .A2(new_n625), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n621), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n612), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n628), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n629), .A2(new_n633), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n620), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G127gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n547), .B1(new_n647), .B2(new_n620), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G183gat), .B(G211gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n653), .B(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n611), .A2(new_n646), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n571), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n372), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND4_X1  g463(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n462), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n462), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n667), .A2(new_n664), .ZN(new_n668));
  OAI221_X1 g467(.A(new_n665), .B1(new_n546), .B2(new_n667), .C1(new_n668), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g468(.A(new_n660), .ZN(new_n670));
  INV_X1    g469(.A(new_n473), .ZN(new_n671));
  OAI21_X1  g470(.A(G15gat), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n456), .A2(G15gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n670), .B2(new_n673), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n660), .A2(new_n474), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n658), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n646), .A2(new_n610), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n571), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n512), .A3(new_n661), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n511), .B2(new_n610), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n375), .A2(new_n474), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n687), .A2(new_n510), .A3(new_n671), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n496), .A2(new_n368), .A3(new_n374), .A4(new_n401), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n689), .A2(KEYINPUT35), .B1(new_n461), .B2(new_n464), .ZN(new_n690));
  OAI211_X1 g489(.A(KEYINPUT44), .B(new_n611), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n646), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n559), .A2(new_n564), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n567), .B1(new_n566), .B2(new_n555), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n565), .A2(KEYINPUT103), .A3(new_n568), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n692), .A2(new_n658), .A3(new_n693), .A4(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n372), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(new_n462), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n681), .A2(G36gat), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT46), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n701), .B2(new_n704), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  OAI21_X1  g507(.A(new_n518), .B1(new_n681), .B2(new_n456), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n473), .A2(G43gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n701), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g511(.A(new_n524), .B1(new_n682), .B2(new_n474), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(KEYINPUT104), .B2(KEYINPUT48), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n474), .A2(new_n524), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n701), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1331gat));
  AOI21_X1  g517(.A(new_n658), .B1(new_n607), .B2(new_n609), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n719), .A3(new_n646), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n511), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n661), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g522(.A(new_n704), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT105), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1333gat));
  INV_X1    g527(.A(new_n721), .ZN(new_n729));
  OAI21_X1  g528(.A(G71gat), .B1(new_n729), .B2(new_n671), .ZN(new_n730));
  INV_X1    g529(.A(G71gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n721), .A2(new_n731), .A3(new_n401), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g533(.A1(new_n721), .A2(new_n474), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT107), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT106), .B(G78gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1335gat));
  NAND2_X1  g537(.A1(new_n699), .A2(new_n658), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n693), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n692), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n372), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NOR4_X1   g543(.A1(new_n511), .A2(new_n744), .A3(new_n610), .A4(new_n739), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT108), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n455), .A2(new_n465), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n687), .A2(new_n510), .A3(new_n671), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n610), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n739), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT51), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n746), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n693), .A2(G85gat), .A3(new_n372), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n758), .ZN(G1336gat));
  NOR3_X1   g558(.A1(new_n693), .A2(G92gat), .A3(new_n704), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT109), .Z(new_n762));
  OAI21_X1  g561(.A(G92gat), .B1(new_n742), .B2(new_n704), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n745), .B2(new_n751), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n762), .A2(new_n765), .B1(new_n767), .B2(new_n764), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n742), .B2(new_n671), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n693), .A2(G99gat), .A3(new_n456), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n756), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1338gat));
  NAND4_X1  g571(.A1(new_n686), .A2(new_n474), .A3(new_n691), .A4(new_n740), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G106gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT110), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n776), .A3(G106gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n693), .A2(G106gat), .A3(new_n496), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n745), .B2(new_n751), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT111), .B(new_n778), .C1(new_n745), .C2(new_n751), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n775), .A2(new_n777), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT53), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n756), .B2(new_n778), .ZN(new_n785));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n773), .B2(KEYINPUT112), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT112), .B2(new_n773), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n784), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1339gat));
  NAND3_X1  g593(.A1(new_n699), .A2(new_n693), .A3(new_n719), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n699), .A2(new_n693), .A3(KEYINPUT114), .A4(new_n719), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n633), .B1(new_n627), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n624), .A2(new_n626), .A3(new_n613), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n640), .A2(new_n802), .A3(KEYINPUT54), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n804), .A2(KEYINPUT55), .B1(new_n634), .B2(new_n643), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n803), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n805), .A2(new_n697), .A3(new_n698), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n549), .B1(new_n548), .B2(new_n551), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n556), .A2(new_n557), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n563), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n568), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n646), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n611), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n611), .A2(new_n813), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT55), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n644), .A2(new_n808), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n658), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n454), .A2(new_n372), .A3(new_n462), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n570), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n699), .A2(G113gat), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n824), .B2(new_n827), .ZN(G1340gat));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n646), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n678), .ZN(new_n831));
  INV_X1    g630(.A(G127gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n831), .B(new_n833), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n823), .A2(new_n611), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n835), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT56), .B1(new_n835), .B2(G134gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(G134gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(G1343gat));
  NAND2_X1  g638(.A1(new_n293), .A2(new_n295), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n473), .A2(new_n372), .A3(new_n462), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n821), .B2(new_n474), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n474), .A2(KEYINPUT57), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n805), .A2(new_n569), .A3(new_n808), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n611), .B1(new_n844), .B2(new_n814), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n658), .B1(new_n845), .B2(new_n819), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n799), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n841), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n840), .B1(new_n848), .B2(new_n570), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n797), .A2(new_n798), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n814), .B1(new_n699), .B2(new_n818), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n610), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n816), .A2(new_n818), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n851), .B1(new_n855), .B2(new_n658), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n496), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n841), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n569), .A2(new_n292), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT117), .Z(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n849), .A2(new_n850), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n840), .B1(new_n848), .B2(new_n699), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n850), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n659), .A2(new_n570), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n496), .B1(new_n867), .B2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n846), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n843), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n646), .B(new_n841), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n858), .B2(new_n646), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n646), .A2(new_n875), .ZN(new_n877));
  OAI221_X1 g676(.A(new_n874), .B1(G148gat), .B2(new_n876), .C1(new_n848), .C2(new_n877), .ZN(G1345gat));
  OAI21_X1  g677(.A(G155gat), .B1(new_n848), .B2(new_n658), .ZN(new_n879));
  INV_X1    g678(.A(G155gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n880), .A3(new_n678), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT119), .Z(G1346gat));
  NOR4_X1   g682(.A1(new_n610), .A2(G162gat), .A3(new_n372), .A4(new_n462), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n671), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT120), .ZN(new_n886));
  OAI21_X1  g685(.A(G162gat), .B1(new_n848), .B2(new_n610), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1347gat));
  AOI21_X1  g687(.A(new_n661), .B1(new_n799), .B2(new_n820), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n462), .B1(new_n889), .B2(KEYINPUT121), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n891), .B(new_n661), .C1(new_n799), .C2(new_n820), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n890), .A2(new_n454), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n700), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n704), .A2(new_n661), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(KEYINPUT122), .A3(new_n401), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT122), .B1(new_n895), .B2(new_n401), .ZN(new_n897));
  OR4_X1    g696(.A1(new_n474), .A2(new_n856), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G169gat), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n570), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n894), .A2(new_n900), .ZN(G1348gat));
  OAI21_X1  g700(.A(G176gat), .B1(new_n898), .B2(new_n693), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n891), .B1(new_n856), .B2(new_n661), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n462), .A4(new_n461), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n693), .A2(G176gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1349gat));
  OAI21_X1  g706(.A(G183gat), .B1(new_n898), .B2(new_n658), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n658), .A2(new_n246), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT123), .B1(new_n893), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  INV_X1    g710(.A(new_n909), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n905), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(new_n908), .C1(new_n910), .C2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n898), .B2(new_n610), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n893), .A2(new_n248), .A3(new_n611), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n890), .A2(new_n892), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n473), .A2(new_n496), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n700), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G197gat), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n871), .A2(new_n872), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n671), .A2(new_n895), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT125), .Z(new_n933));
  AND2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n570), .A2(new_n930), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n929), .A2(new_n930), .B1(new_n934), .B2(new_n935), .ZN(G1352gat));
  INV_X1    g735(.A(G204gat), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n646), .B(new_n933), .C1(new_n871), .C2(new_n872), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(KEYINPUT127), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(KEYINPUT127), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g739(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n693), .A2(G204gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n923), .A2(new_n924), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n944));
  INV_X1    g743(.A(new_n942), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n925), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n943), .A3(new_n946), .ZN(G1353gat));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n928), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n678), .A2(new_n204), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n678), .B(new_n933), .C1(new_n871), .C2(new_n872), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n948), .A2(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n611), .A3(new_n933), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G218gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n611), .A2(new_n205), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n948), .B2(new_n956), .ZN(G1355gat));
endmodule


