

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U550 ( .A(n881), .Z(n516) );
  NOR2_X1 U551 ( .A1(n764), .A2(n766), .ZN(n692) );
  NOR2_X4 U552 ( .A1(G2105), .A2(n520), .ZN(n883) );
  XOR2_X1 U553 ( .A(KEYINPUT17), .B(n517), .Z(n881) );
  NOR2_X1 U554 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  OR2_X1 U555 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U556 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U557 ( .A1(n697), .A2(n991), .ZN(n704) );
  NOR2_X1 U558 ( .A1(G2084), .A2(n699), .ZN(n679) );
  NOR2_X1 U559 ( .A1(G164), .A2(G1384), .ZN(n676) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  NOR2_X1 U561 ( .A1(n768), .A2(n767), .ZN(n801) );
  NOR2_X1 U562 ( .A1(G651), .A2(n631), .ZN(n639) );
  NOR2_X1 U563 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U564 ( .A(G2104), .ZN(n520) );
  NAND2_X1 U565 ( .A1(G102), .A2(n883), .ZN(n519) );
  NAND2_X1 U566 ( .A1(G138), .A2(n881), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n525) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U569 ( .A1(G114), .A2(n890), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n520), .A2(G2105), .ZN(n521) );
  XNOR2_X1 U571 ( .A(n521), .B(KEYINPUT65), .ZN(n535) );
  NAND2_X1 U572 ( .A1(G126), .A2(n535), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U574 ( .A1(n525), .A2(n524), .ZN(G164) );
  NAND2_X1 U575 ( .A1(n890), .A2(G113), .ZN(n528) );
  NAND2_X1 U576 ( .A1(G101), .A2(n883), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(n526), .Z(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U579 ( .A1(G137), .A2(n516), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G125), .A2(n535), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n531) );
  AND2_X1 U582 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U583 ( .A1(G99), .A2(n883), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G111), .A2(n890), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n541) );
  BUF_X1 U586 ( .A(n535), .Z(n887) );
  NAND2_X1 U587 ( .A1(G123), .A2(n887), .ZN(n536) );
  XNOR2_X1 U588 ( .A(n536), .B(KEYINPUT18), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT74), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G135), .A2(n516), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n912) );
  XNOR2_X1 U593 ( .A(n912), .B(G2096), .ZN(n542) );
  XNOR2_X1 U594 ( .A(n542), .B(KEYINPUT75), .ZN(n543) );
  OR2_X1 U595 ( .A1(G2100), .A2(n543), .ZN(G156) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G57), .ZN(G237) );
  INV_X1 U598 ( .A(G120), .ZN(G236) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n631) );
  NAND2_X1 U600 ( .A1(G53), .A2(n639), .ZN(n546) );
  INV_X1 U601 ( .A(G651), .ZN(n547) );
  NOR2_X1 U602 ( .A1(G543), .A2(n547), .ZN(n544) );
  XOR2_X1 U603 ( .A(KEYINPUT1), .B(n544), .Z(n643) );
  NAND2_X1 U604 ( .A1(G65), .A2(n643), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n551) );
  NOR2_X1 U606 ( .A1(G543), .A2(G651), .ZN(n634) );
  NAND2_X1 U607 ( .A1(G91), .A2(n634), .ZN(n549) );
  NOR2_X1 U608 ( .A1(n631), .A2(n547), .ZN(n635) );
  NAND2_X1 U609 ( .A1(G78), .A2(n635), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n714) );
  INV_X1 U612 ( .A(n714), .ZN(G299) );
  XNOR2_X1 U613 ( .A(KEYINPUT71), .B(KEYINPUT5), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n634), .A2(G89), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G76), .A2(n635), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n556), .B(n555), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n639), .A2(G51), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT72), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G63), .A2(n643), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT73), .B(n560), .Z(n561) );
  XNOR2_X1 U624 ( .A(KEYINPUT6), .B(n561), .ZN(n562) );
  NOR2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT7), .B(n564), .Z(G168) );
  NAND2_X1 U627 ( .A1(G90), .A2(n634), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G77), .A2(n635), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n567), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n639), .A2(G52), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G64), .A2(n643), .ZN(n568) );
  AND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(G301) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U636 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n573) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n817) );
  NAND2_X1 U640 ( .A1(n817), .A2(G567), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U642 ( .A1(G56), .A2(n643), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n575), .Z(n581) );
  NAND2_X1 U644 ( .A1(n634), .A2(G81), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G68), .A2(n635), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n639), .A2(G43), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n991) );
  INV_X1 U652 ( .A(G860), .ZN(n597) );
  OR2_X1 U653 ( .A1(n991), .A2(n597), .ZN(G153) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G66), .A2(n643), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G92), .A2(n634), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G54), .A2(n639), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n635), .A2(G79), .ZN(n586) );
  XOR2_X1 U660 ( .A(KEYINPUT70), .B(n586), .Z(n587) );
  NOR2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT15), .ZN(n998) );
  OR2_X1 U664 ( .A1(n998), .A2(G868), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(G284) );
  INV_X1 U666 ( .A(G868), .ZN(n594) );
  NOR2_X1 U667 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n597), .A2(G559), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n598), .A2(n998), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n991), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n998), .A2(G868), .ZN(n600) );
  NOR2_X1 U675 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U677 ( .A1(n998), .A2(G559), .ZN(n656) );
  XNOR2_X1 U678 ( .A(n991), .B(n656), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n603), .A2(G860), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G55), .A2(n639), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G67), .A2(n643), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(KEYINPUT76), .B(n606), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G93), .A2(n634), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G80), .A2(n635), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n653) );
  XNOR2_X1 U688 ( .A(n611), .B(n653), .ZN(G145) );
  NAND2_X1 U689 ( .A1(G86), .A2(n634), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G61), .A2(n643), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT77), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G48), .A2(n639), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n635), .A2(G73), .ZN(n617) );
  XOR2_X1 U696 ( .A(KEYINPUT2), .B(n617), .Z(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT78), .B(n620), .Z(G305) );
  NAND2_X1 U699 ( .A1(G88), .A2(n634), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G62), .A2(n643), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G75), .A2(n635), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n623), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n639), .A2(G50), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(G303) );
  INV_X1 U707 ( .A(G303), .ZN(G166) );
  NAND2_X1 U708 ( .A1(G49), .A2(n639), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n643), .A2(n630), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G85), .A2(n634), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G72), .A2(n635), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U717 ( .A(KEYINPUT66), .B(n638), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G47), .A2(n639), .ZN(n640) );
  XNOR2_X1 U719 ( .A(KEYINPUT67), .B(n640), .ZN(n641) );
  NOR2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n643), .A2(G60), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G290) );
  NOR2_X1 U723 ( .A1(G868), .A2(n653), .ZN(n646) );
  XOR2_X1 U724 ( .A(n646), .B(KEYINPUT82), .Z(n659) );
  XNOR2_X1 U725 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n648) );
  XNOR2_X1 U726 ( .A(G288), .B(KEYINPUT80), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(G166), .B(n649), .ZN(n651) );
  XNOR2_X1 U729 ( .A(G290), .B(n714), .ZN(n650) );
  XNOR2_X1 U730 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(n991), .ZN(n655) );
  XNOR2_X1 U733 ( .A(G305), .B(n655), .ZN(n898) );
  XOR2_X1 U734 ( .A(n898), .B(n656), .Z(n657) );
  NAND2_X1 U735 ( .A1(G868), .A2(n657), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U743 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NOR2_X1 U744 ( .A1(G236), .A2(G237), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G69), .A2(n664), .ZN(n665) );
  XNOR2_X1 U746 ( .A(KEYINPUT83), .B(n665), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n666), .A2(G108), .ZN(n821) );
  NAND2_X1 U748 ( .A1(n821), .A2(G567), .ZN(n671) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U751 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U752 ( .A1(G96), .A2(n669), .ZN(n822) );
  NAND2_X1 U753 ( .A1(n822), .A2(G2106), .ZN(n670) );
  NAND2_X1 U754 ( .A1(n671), .A2(n670), .ZN(n908) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n672) );
  XNOR2_X1 U756 ( .A(KEYINPUT84), .B(n672), .ZN(n673) );
  NOR2_X1 U757 ( .A1(n908), .A2(n673), .ZN(n820) );
  NAND2_X1 U758 ( .A1(G36), .A2(n820), .ZN(n674) );
  XOR2_X1 U759 ( .A(KEYINPUT85), .B(n674), .Z(G176) );
  XOR2_X1 U760 ( .A(G2078), .B(KEYINPUT25), .Z(n964) );
  INV_X1 U761 ( .A(KEYINPUT64), .ZN(n675) );
  XNOR2_X1 U762 ( .A(n676), .B(n675), .ZN(n764) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n766) );
  INV_X1 U764 ( .A(n692), .ZN(n699) );
  NOR2_X1 U765 ( .A1(n964), .A2(n699), .ZN(n678) );
  BUF_X1 U766 ( .A(n692), .Z(n708) );
  NOR2_X1 U767 ( .A1(n708), .A2(G1961), .ZN(n677) );
  NOR2_X1 U768 ( .A1(n678), .A2(n677), .ZN(n720) );
  NAND2_X1 U769 ( .A1(G301), .A2(n720), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G8), .A2(n699), .ZN(n759) );
  NOR2_X1 U771 ( .A1(G1966), .A2(n759), .ZN(n737) );
  XOR2_X1 U772 ( .A(KEYINPUT92), .B(n679), .Z(n731) );
  NAND2_X1 U773 ( .A1(G8), .A2(n731), .ZN(n680) );
  NOR2_X1 U774 ( .A1(n737), .A2(n680), .ZN(n682) );
  XNOR2_X1 U775 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n681) );
  XNOR2_X1 U776 ( .A(n682), .B(n681), .ZN(n683) );
  OR2_X1 U777 ( .A1(G168), .A2(n683), .ZN(n684) );
  XOR2_X1 U778 ( .A(KEYINPUT31), .B(n686), .Z(n734) );
  INV_X1 U779 ( .A(G8), .ZN(n691) );
  NOR2_X1 U780 ( .A1(G1971), .A2(n759), .ZN(n688) );
  NOR2_X1 U781 ( .A1(G2090), .A2(n699), .ZN(n687) );
  NOR2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n689), .A2(G303), .ZN(n690) );
  OR2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n725) );
  AND2_X1 U785 ( .A1(n734), .A2(n725), .ZN(n724) );
  NAND2_X1 U786 ( .A1(G1996), .A2(n692), .ZN(n693) );
  XNOR2_X1 U787 ( .A(n693), .B(KEYINPUT26), .ZN(n695) );
  NAND2_X1 U788 ( .A1(G1341), .A2(n699), .ZN(n694) );
  NAND2_X1 U789 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U790 ( .A(n696), .B(KEYINPUT96), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n998), .A2(n704), .ZN(n703) );
  AND2_X1 U792 ( .A1(n708), .A2(G2067), .ZN(n698) );
  XNOR2_X1 U793 ( .A(n698), .B(KEYINPUT97), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n699), .A2(G1348), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n706) );
  OR2_X1 U797 ( .A1(n704), .A2(n998), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n712) );
  NAND2_X1 U799 ( .A1(n708), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT27), .ZN(n710) );
  XOR2_X1 U801 ( .A(G1956), .B(KEYINPUT94), .Z(n936) );
  NOR2_X1 U802 ( .A1(n708), .A2(n936), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U807 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n715) );
  XNOR2_X1 U808 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U810 ( .A(n719), .B(KEYINPUT29), .ZN(n722) );
  NOR2_X1 U811 ( .A1(G301), .A2(n720), .ZN(n721) );
  XNOR2_X1 U812 ( .A(n723), .B(KEYINPUT98), .ZN(n735) );
  NAND2_X1 U813 ( .A1(n724), .A2(n735), .ZN(n729) );
  INV_X1 U814 ( .A(n725), .ZN(n727) );
  AND2_X1 U815 ( .A1(G286), .A2(G8), .ZN(n726) );
  OR2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U818 ( .A(n730), .B(KEYINPUT32), .ZN(n741) );
  INV_X1 U819 ( .A(n731), .ZN(n732) );
  NAND2_X1 U820 ( .A1(G8), .A2(n732), .ZN(n733) );
  XOR2_X1 U821 ( .A(KEYINPUT93), .B(n733), .Z(n739) );
  AND2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n741), .A2(n740), .ZN(n753) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n747) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U828 ( .A1(n747), .A2(n742), .ZN(n996) );
  NAND2_X1 U829 ( .A1(n753), .A2(n996), .ZN(n743) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NAND2_X1 U831 ( .A1(n743), .A2(n993), .ZN(n744) );
  INV_X1 U832 ( .A(n759), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n745), .A2(n746), .ZN(n750) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT100), .ZN(n752) );
  XOR2_X1 U838 ( .A(G305), .B(G1981), .Z(n1009) );
  AND2_X1 U839 ( .A1(n752), .A2(n1009), .ZN(n763) );
  NOR2_X1 U840 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n753), .A2(n755), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n756), .A2(n759), .ZN(n761) );
  NOR2_X1 U844 ( .A1(G305), .A2(G1981), .ZN(n757) );
  XOR2_X1 U845 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  OR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n768) );
  XNOR2_X1 U849 ( .A(G1986), .B(G290), .ZN(n1004) );
  INV_X1 U850 ( .A(n764), .ZN(n765) );
  NOR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n812) );
  AND2_X1 U852 ( .A1(n1004), .A2(n812), .ZN(n767) );
  XNOR2_X1 U853 ( .A(KEYINPUT34), .B(KEYINPUT86), .ZN(n772) );
  NAND2_X1 U854 ( .A1(G104), .A2(n883), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G140), .A2(n516), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n772), .B(n771), .ZN(n778) );
  NAND2_X1 U858 ( .A1(n890), .A2(G116), .ZN(n773) );
  XOR2_X1 U859 ( .A(KEYINPUT87), .B(n773), .Z(n775) );
  NAND2_X1 U860 ( .A1(n887), .A2(G128), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n779), .B(KEYINPUT36), .ZN(n780) );
  XNOR2_X1 U865 ( .A(n780), .B(KEYINPUT88), .ZN(n870) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U867 ( .A1(n870), .A2(n810), .ZN(n931) );
  NAND2_X1 U868 ( .A1(n812), .A2(n931), .ZN(n807) );
  INV_X1 U869 ( .A(n807), .ZN(n798) );
  NAND2_X1 U870 ( .A1(G95), .A2(n883), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G107), .A2(n890), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G131), .A2(n516), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G119), .A2(n887), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n878) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n878), .ZN(n796) );
  NAND2_X1 U878 ( .A1(G105), .A2(n883), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT38), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G117), .A2(n890), .ZN(n789) );
  NAND2_X1 U881 ( .A1(G141), .A2(n516), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G129), .A2(n887), .ZN(n790) );
  XNOR2_X1 U884 ( .A(KEYINPUT89), .B(n790), .ZN(n791) );
  NOR2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n862) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n862), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n917) );
  NAND2_X1 U889 ( .A1(n917), .A2(n812), .ZN(n797) );
  XOR2_X1 U890 ( .A(KEYINPUT90), .B(n797), .Z(n804) );
  NOR2_X1 U891 ( .A1(n798), .A2(n804), .ZN(n799) );
  XOR2_X1 U892 ( .A(n799), .B(KEYINPUT91), .Z(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n815) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n862), .ZN(n910) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U896 ( .A1(G1991), .A2(n878), .ZN(n913) );
  NOR2_X1 U897 ( .A1(n802), .A2(n913), .ZN(n803) );
  NOR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n910), .A2(n805), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(KEYINPUT39), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U902 ( .A(KEYINPUT101), .B(n809), .Z(n811) );
  NAND2_X1 U903 ( .A1(n870), .A2(n810), .ZN(n918) );
  NAND2_X1 U904 ( .A1(n811), .A2(n918), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U907 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(G188) );
  INV_X1 U914 ( .A(G108), .ZN(G238) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  NOR2_X1 U916 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  XOR2_X1 U918 ( .A(KEYINPUT43), .B(G2678), .Z(n824) );
  XNOR2_X1 U919 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT42), .B(G2090), .Z(n826) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2072), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U924 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U925 ( .A(G2096), .B(G2100), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(n832) );
  XOR2_X1 U927 ( .A(G2084), .B(G2078), .Z(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(G227) );
  XOR2_X1 U929 ( .A(G1981), .B(G1961), .Z(n834) );
  XNOR2_X1 U930 ( .A(G1991), .B(G1966), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(G1976), .B(G1971), .Z(n836) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1956), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT105), .B(G2474), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U938 ( .A(G1996), .B(KEYINPUT41), .Z(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(G229) );
  XNOR2_X1 U940 ( .A(G1341), .B(G2454), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n843), .B(G2430), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n844), .B(G1348), .ZN(n850) );
  XOR2_X1 U943 ( .A(G2443), .B(G2427), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2438), .B(G2446), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U946 ( .A(G2451), .B(G2435), .Z(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n851), .A2(G14), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT102), .B(n852), .Z(G401) );
  NAND2_X1 U951 ( .A1(G100), .A2(n883), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G112), .A2(n890), .ZN(n853) );
  NAND2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G124), .A2(n887), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT106), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G136), .A2(n516), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U959 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U960 ( .A(G162), .B(n912), .Z(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n874) );
  NAND2_X1 U962 ( .A1(G103), .A2(n883), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G139), .A2(n516), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G115), .A2(n890), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G127), .A2(n887), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT47), .B(n867), .Z(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n920) );
  XOR2_X1 U970 ( .A(n920), .B(n870), .Z(n872) );
  XNOR2_X1 U971 ( .A(G160), .B(G164), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n880) );
  XOR2_X1 U974 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n895) );
  NAND2_X1 U979 ( .A1(n516), .A2(G142), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n882), .B(KEYINPUT108), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n886), .B(KEYINPUT45), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n893) );
  NAND2_X1 U986 ( .A1(G118), .A2(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(KEYINPUT107), .B(n891), .ZN(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G395) );
  INV_X1 U991 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U992 ( .A(G171), .B(n998), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n897), .B(G286), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(G397) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n902) );
  XNOR2_X1 U997 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n905) );
  NOR2_X1 U999 ( .A1(n908), .A2(G401), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(KEYINPUT111), .B(n903), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(n908), .ZN(G319) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1007 ( .A(G2090), .B(G162), .Z(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT51), .B(n911), .Z(n929) );
  XNOR2_X1 U1010 ( .A(G160), .B(G2084), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n927) );
  XNOR2_X1 U1015 ( .A(G164), .B(G2078), .ZN(n923) );
  XOR2_X1 U1016 ( .A(G2072), .B(n920), .Z(n921) );
  XNOR2_X1 U1017 ( .A(KEYINPUT113), .B(n921), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n924), .B(KEYINPUT114), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n925), .B(KEYINPUT50), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1022 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1024 ( .A(KEYINPUT52), .B(n932), .Z(n933) );
  NOR2_X1 U1025 ( .A1(KEYINPUT55), .A2(n933), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(KEYINPUT115), .B(n934), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(n935), .A2(G29), .ZN(n990) );
  XOR2_X1 U1028 ( .A(G1961), .B(G5), .Z(n951) );
  XNOR2_X1 U1029 ( .A(n936), .B(G20), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(n937), .B(KEYINPUT124), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(G1348), .B(KEYINPUT59), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n938), .B(G4), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n945) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n942) );
  XNOR2_X1 U1035 ( .A(G6), .B(G1981), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT125), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1039 ( .A(KEYINPUT60), .B(n946), .Z(n948) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT126), .B(n949), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n959) );
  XNOR2_X1 U1044 ( .A(G1986), .B(G24), .ZN(n956) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G1976), .B(G23), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT58), .B(n957), .Z(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1052 ( .A(KEYINPUT61), .B(n960), .Z(n961) );
  NOR2_X1 U1053 ( .A1(G16), .A2(n961), .ZN(n988) );
  XOR2_X1 U1054 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n983) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G35), .ZN(n978) );
  XNOR2_X1 U1056 ( .A(KEYINPUT119), .B(G1996), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(G32), .ZN(n969) );
  XOR2_X1 U1058 ( .A(G1991), .B(G25), .Z(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G27), .B(n964), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT118), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G2072), .B(KEYINPUT116), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(G33), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G26), .B(G2067), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n973), .B(KEYINPUT117), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT53), .B(n976), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1072 ( .A(G2084), .B(G34), .Z(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT54), .B(n979), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n985) );
  INV_X1 U1076 ( .A(G29), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(G11), .A2(n986), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n1018) );
  XOR2_X1 U1081 ( .A(KEYINPUT56), .B(G16), .Z(n1016) );
  XOR2_X1 U1082 ( .A(n991), .B(G1341), .Z(n1007) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G299), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G171), .B(G1961), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(G1348), .B(n998), .Z(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(KEYINPUT122), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1095 ( .A(G1966), .B(G168), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT121), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT57), .B(n1011), .Z(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(KEYINPUT123), .B(n1014), .Z(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

