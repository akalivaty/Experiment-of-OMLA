

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(n735), .ZN(n712) );
  AND2_X2 U554 ( .A1(n537), .A2(G2104), .ZN(n883) );
  NOR2_X1 U555 ( .A1(n689), .A2(n946), .ZN(n690) );
  NOR2_X1 U556 ( .A1(n724), .A2(n723), .ZN(n725) );
  INV_X1 U557 ( .A(KEYINPUT98), .ZN(n682) );
  INV_X1 U558 ( .A(KEYINPUT102), .ZN(n728) );
  XNOR2_X1 U559 ( .A(n683), .B(n682), .ZN(n717) );
  XNOR2_X1 U560 ( .A(n732), .B(n728), .ZN(n729) );
  XNOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT32), .ZN(n742) );
  XNOR2_X1 U562 ( .A(n743), .B(n742), .ZN(n744) );
  AND2_X1 U563 ( .A1(G160), .A2(G40), .ZN(n785) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n537), .ZN(n875) );
  NOR2_X1 U565 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U566 ( .A1(n643), .A2(G89), .ZN(n520) );
  XNOR2_X1 U567 ( .A(n520), .B(KEYINPUT4), .ZN(n522) );
  XOR2_X1 U568 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  INV_X1 U569 ( .A(G651), .ZN(n524) );
  NOR2_X1 U570 ( .A1(n638), .A2(n524), .ZN(n644) );
  NAND2_X1 U571 ( .A1(G76), .A2(n644), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT5), .ZN(n531) );
  NOR2_X1 U574 ( .A1(n524), .A2(G543), .ZN(n525) );
  XOR2_X2 U575 ( .A(KEYINPUT1), .B(n525), .Z(n648) );
  NAND2_X1 U576 ( .A1(G63), .A2(n648), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G651), .A2(n638), .ZN(n526) );
  XOR2_X1 U578 ( .A(KEYINPUT65), .B(n526), .Z(n649) );
  NAND2_X1 U579 ( .A1(G51), .A2(n649), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U583 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U584 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XOR2_X2 U586 ( .A(KEYINPUT17), .B(n533), .Z(n880) );
  NAND2_X1 U587 ( .A1(n880), .A2(G137), .ZN(n536) );
  INV_X1 U588 ( .A(G2105), .ZN(n537) );
  NAND2_X1 U589 ( .A1(G101), .A2(n883), .ZN(n534) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(n534), .Z(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G125), .A2(n875), .ZN(n539) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U594 ( .A1(G113), .A2(n876), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U596 ( .A1(n541), .A2(n540), .ZN(G160) );
  NAND2_X1 U597 ( .A1(n880), .A2(G138), .ZN(n548) );
  NAND2_X1 U598 ( .A1(G102), .A2(n883), .ZN(n542) );
  XNOR2_X1 U599 ( .A(KEYINPUT89), .B(n542), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G126), .A2(n875), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G114), .A2(n876), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G64), .A2(n648), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G52), .A2(n649), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U608 ( .A(KEYINPUT67), .B(n551), .Z(n556) );
  NAND2_X1 U609 ( .A1(G90), .A2(n643), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G77), .A2(n644), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G120), .ZN(G236) );
  INV_X1 U616 ( .A(G69), .ZN(G235) );
  INV_X1 U617 ( .A(G108), .ZN(G238) );
  INV_X1 U618 ( .A(G132), .ZN(G219) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  NAND2_X1 U620 ( .A1(G88), .A2(n643), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G75), .A2(n644), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G62), .A2(n648), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G50), .A2(n649), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(G166) );
  XOR2_X1 U627 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n564) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT70), .B(n565), .ZN(G223) );
  XOR2_X1 U631 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n567) );
  INV_X1 U632 ( .A(G223), .ZN(n830) );
  NAND2_X1 U633 ( .A1(n830), .A2(G567), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G234) );
  NAND2_X1 U635 ( .A1(G56), .A2(n648), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n568), .Z(n575) );
  NAND2_X1 U637 ( .A1(G81), .A2(n643), .ZN(n569) );
  XOR2_X1 U638 ( .A(KEYINPUT12), .B(n569), .Z(n570) );
  XNOR2_X1 U639 ( .A(n570), .B(KEYINPUT73), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G68), .A2(n644), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  NOR2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n649), .A2(G43), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n946) );
  INV_X1 U646 ( .A(G860), .ZN(n618) );
  OR2_X1 U647 ( .A1(n946), .A2(n618), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G54), .A2(n649), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G92), .A2(n643), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G79), .A2(n644), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n648), .A2(G66), .ZN(n580) );
  XOR2_X1 U655 ( .A(KEYINPUT74), .B(n580), .Z(n581) );
  NOR2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT15), .ZN(n586) );
  XOR2_X2 U659 ( .A(KEYINPUT75), .B(n586), .Z(n945) );
  INV_X1 U660 ( .A(n945), .ZN(n696) );
  INV_X1 U661 ( .A(G868), .ZN(n662) );
  NAND2_X1 U662 ( .A1(n696), .A2(n662), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n643), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G78), .A2(n644), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U667 ( .A(KEYINPUT68), .B(n591), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n649), .A2(G53), .ZN(n592) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n592), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n648), .A2(G65), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U674 ( .A1(G286), .A2(n662), .ZN(n597) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n618), .A2(G559), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n599), .A2(n945), .ZN(n600) );
  XNOR2_X1 U678 ( .A(n600), .B(KEYINPUT76), .ZN(n601) );
  XNOR2_X1 U679 ( .A(KEYINPUT16), .B(n601), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n946), .ZN(n602) );
  XOR2_X1 U681 ( .A(KEYINPUT77), .B(n602), .Z(n605) );
  NAND2_X1 U682 ( .A1(G868), .A2(n945), .ZN(n603) );
  NOR2_X1 U683 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(G282) );
  XNOR2_X1 U685 ( .A(G2100), .B(KEYINPUT79), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n875), .A2(G123), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n606), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G135), .A2(n880), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U690 ( .A(KEYINPUT78), .B(n609), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G99), .A2(n883), .ZN(n611) );
  NAND2_X1 U692 ( .A1(G111), .A2(n876), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n972) );
  XNOR2_X1 U695 ( .A(n972), .B(G2096), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U697 ( .A(KEYINPUT80), .B(n616), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G559), .A2(n945), .ZN(n617) );
  XOR2_X1 U699 ( .A(n946), .B(n617), .Z(n660) );
  NAND2_X1 U700 ( .A1(n618), .A2(n660), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G80), .A2(n644), .ZN(n620) );
  NAND2_X1 U702 ( .A1(G67), .A2(n648), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U704 ( .A1(G93), .A2(n643), .ZN(n621) );
  XNOR2_X1 U705 ( .A(KEYINPUT81), .B(n621), .ZN(n622) );
  NOR2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n649), .A2(G55), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n663) );
  XNOR2_X1 U709 ( .A(n626), .B(n663), .ZN(G145) );
  NAND2_X1 U710 ( .A1(G48), .A2(n649), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G86), .A2(n643), .ZN(n628) );
  NAND2_X1 U712 ( .A1(G61), .A2(n648), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n644), .A2(G73), .ZN(n629) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U716 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n634), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U719 ( .A1(G49), .A2(n649), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U722 ( .A(KEYINPUT82), .B(n637), .Z(n642) );
  NAND2_X1 U723 ( .A1(G87), .A2(n638), .ZN(n639) );
  XNOR2_X1 U724 ( .A(KEYINPUT83), .B(n639), .ZN(n640) );
  NOR2_X1 U725 ( .A1(n648), .A2(n640), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G85), .A2(n643), .ZN(n646) );
  NAND2_X1 U728 ( .A1(G72), .A2(n644), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U730 ( .A(KEYINPUT66), .B(n647), .Z(n653) );
  NAND2_X1 U731 ( .A1(G60), .A2(n648), .ZN(n651) );
  NAND2_X1 U732 ( .A1(G47), .A2(n649), .ZN(n650) );
  AND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(G290) );
  XNOR2_X1 U735 ( .A(G305), .B(G288), .ZN(n659) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n655) );
  INV_X1 U737 ( .A(G299), .ZN(n707) );
  XNOR2_X1 U738 ( .A(n707), .B(G166), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U740 ( .A(n656), .B(G290), .Z(n657) );
  XNOR2_X1 U741 ( .A(n663), .B(n657), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n659), .B(n658), .ZN(n898) );
  XOR2_X1 U743 ( .A(n898), .B(n660), .Z(n661) );
  NOR2_X1 U744 ( .A1(n662), .A2(n661), .ZN(n665) );
  NOR2_X1 U745 ( .A1(G868), .A2(n663), .ZN(n664) );
  NOR2_X1 U746 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n666) );
  XNOR2_X1 U749 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U756 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G96), .A2(n673), .ZN(n834) );
  NAND2_X1 U758 ( .A1(n834), .A2(G2106), .ZN(n679) );
  NOR2_X1 U759 ( .A1(G235), .A2(G236), .ZN(n674) );
  XNOR2_X1 U760 ( .A(n674), .B(KEYINPUT87), .ZN(n675) );
  NOR2_X1 U761 ( .A1(G238), .A2(n675), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n676), .A2(G57), .ZN(n677) );
  XNOR2_X1 U763 ( .A(n677), .B(KEYINPUT88), .ZN(n835) );
  NAND2_X1 U764 ( .A1(n835), .A2(G567), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n836) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U767 ( .A1(n836), .A2(n680), .ZN(n833) );
  NAND2_X1 U768 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  NOR2_X2 U770 ( .A1(G164), .A2(G1384), .ZN(n787) );
  NAND2_X1 U771 ( .A1(n785), .A2(n787), .ZN(n735) );
  NAND2_X1 U772 ( .A1(G8), .A2(n735), .ZN(n765) );
  NOR2_X1 U773 ( .A1(G1966), .A2(n765), .ZN(n683) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n735), .ZN(n719) );
  NAND2_X1 U775 ( .A1(G8), .A2(n719), .ZN(n684) );
  NAND2_X1 U776 ( .A1(n717), .A2(n684), .ZN(n730) );
  AND2_X1 U777 ( .A1(n712), .A2(G1996), .ZN(n686) );
  XOR2_X1 U778 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n685) );
  XNOR2_X1 U779 ( .A(n686), .B(n685), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n735), .A2(G1341), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U782 ( .A(n690), .B(KEYINPUT64), .Z(n697) );
  OR2_X1 U783 ( .A1(n697), .A2(n696), .ZN(n695) );
  AND2_X1 U784 ( .A1(n735), .A2(G1348), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n691), .B(KEYINPUT101), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n712), .A2(G2067), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n712), .ZN(n700) );
  XOR2_X1 U792 ( .A(KEYINPUT99), .B(n700), .Z(n701) );
  XNOR2_X1 U793 ( .A(KEYINPUT27), .B(n701), .ZN(n703) );
  AND2_X1 U794 ( .A1(n735), .A2(G1956), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U799 ( .A(n708), .B(KEYINPUT28), .Z(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U801 ( .A(KEYINPUT29), .B(n711), .Z(n716) );
  INV_X1 U802 ( .A(G1961), .ZN(n1014) );
  NAND2_X1 U803 ( .A1(n735), .A2(n1014), .ZN(n714) );
  XNOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .ZN(n927) );
  NAND2_X1 U805 ( .A1(n712), .A2(n927), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n722) );
  NAND2_X1 U807 ( .A1(n722), .A2(G171), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n717), .A2(G8), .ZN(n718) );
  NOR2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U811 ( .A(KEYINPUT30), .B(n720), .Z(n721) );
  NOR2_X1 U812 ( .A1(G168), .A2(n721), .ZN(n724) );
  NOR2_X1 U813 ( .A1(G171), .A2(n722), .ZN(n723) );
  XOR2_X1 U814 ( .A(KEYINPUT31), .B(n725), .Z(n726) );
  NAND2_X1 U815 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U817 ( .A(n731), .B(KEYINPUT103), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n732), .A2(G286), .ZN(n740) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n765), .ZN(n733) );
  XOR2_X1 U820 ( .A(KEYINPUT104), .B(n733), .Z(n734) );
  NAND2_X1 U821 ( .A1(n734), .A2(G303), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U824 ( .A(n738), .B(KEYINPUT105), .ZN(n739) );
  NAND2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n741), .A2(G8), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n745), .A2(n744), .ZN(n767) );
  NOR2_X1 U828 ( .A1(G2090), .A2(G303), .ZN(n746) );
  XNOR2_X1 U829 ( .A(n746), .B(KEYINPUT108), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n747), .A2(G8), .ZN(n748) );
  NAND2_X1 U831 ( .A1(n767), .A2(n748), .ZN(n749) );
  NAND2_X1 U832 ( .A1(n749), .A2(n765), .ZN(n753) );
  NOR2_X1 U833 ( .A1(G1981), .A2(G305), .ZN(n750) );
  XOR2_X1 U834 ( .A(n750), .B(KEYINPUT24), .Z(n751) );
  OR2_X1 U835 ( .A1(n765), .A2(n751), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n753), .A2(n752), .ZN(n762) );
  INV_X1 U837 ( .A(KEYINPUT107), .ZN(n755) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NAND2_X1 U839 ( .A1(n959), .A2(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n959), .A2(KEYINPUT107), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U843 ( .A1(n765), .A2(n758), .ZN(n760) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n942) );
  INV_X1 U845 ( .A(n942), .ZN(n759) );
  NOR2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n769) );
  AND2_X1 U847 ( .A1(n769), .A2(KEYINPUT33), .ZN(n761) );
  OR2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n774) );
  INV_X1 U849 ( .A(G1971), .ZN(n997) );
  AND2_X1 U850 ( .A1(G166), .A2(n997), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n763), .A2(n959), .ZN(n764) );
  OR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n960) );
  NAND2_X1 U855 ( .A1(n768), .A2(n960), .ZN(n772) );
  INV_X1 U856 ( .A(n769), .ZN(n770) );
  OR2_X1 U857 ( .A1(KEYINPUT107), .A2(n770), .ZN(n771) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n812) );
  XNOR2_X1 U860 ( .A(KEYINPUT37), .B(G2067), .ZN(n823) );
  NAND2_X1 U861 ( .A1(G104), .A2(n883), .ZN(n776) );
  NAND2_X1 U862 ( .A1(G140), .A2(n880), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n777), .ZN(n783) );
  NAND2_X1 U865 ( .A1(n875), .A2(G128), .ZN(n778) );
  XOR2_X1 U866 ( .A(KEYINPUT91), .B(n778), .Z(n780) );
  NAND2_X1 U867 ( .A1(n876), .A2(G116), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n784), .ZN(n893) );
  NOR2_X1 U872 ( .A1(n823), .A2(n893), .ZN(n985) );
  INV_X1 U873 ( .A(n785), .ZN(n786) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n826) );
  NAND2_X1 U875 ( .A1(n985), .A2(n826), .ZN(n788) );
  XOR2_X1 U876 ( .A(KEYINPUT92), .B(n788), .Z(n820) );
  XNOR2_X1 U877 ( .A(G1986), .B(G290), .ZN(n955) );
  NAND2_X1 U878 ( .A1(n955), .A2(n826), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT90), .B(n789), .Z(n790) );
  NOR2_X1 U880 ( .A1(n820), .A2(n790), .ZN(n810) );
  NAND2_X1 U881 ( .A1(n876), .A2(G117), .ZN(n791) );
  XNOR2_X1 U882 ( .A(KEYINPUT95), .B(n791), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n875), .A2(G129), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT94), .B(n792), .Z(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U886 ( .A(KEYINPUT96), .B(n795), .Z(n799) );
  NAND2_X1 U887 ( .A1(G105), .A2(n883), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n796), .B(KEYINPUT38), .ZN(n797) );
  XNOR2_X1 U889 ( .A(KEYINPUT97), .B(n797), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n880), .A2(G141), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n892) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n892), .ZN(n809) );
  XOR2_X1 U894 ( .A(KEYINPUT93), .B(G1991), .Z(n922) );
  NAND2_X1 U895 ( .A1(G119), .A2(n875), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G131), .A2(n880), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G95), .A2(n883), .ZN(n805) );
  NAND2_X1 U899 ( .A1(G107), .A2(n876), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  OR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n887) );
  NAND2_X1 U902 ( .A1(n922), .A2(n887), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n973) );
  NAND2_X1 U904 ( .A1(n826), .A2(n973), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n810), .A2(n814), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n813), .B(KEYINPUT109), .ZN(n828) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n892), .ZN(n978) );
  INV_X1 U909 ( .A(n814), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n922), .A2(n887), .ZN(n974) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n974), .A2(n815), .ZN(n816) );
  NOR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n978), .A2(n818), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n819), .B(KEYINPUT39), .ZN(n822) );
  INV_X1 U916 ( .A(n820), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n823), .A2(n893), .ZN(n982) );
  NAND2_X1 U919 ( .A1(n824), .A2(n982), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U925 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  NOR2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  INV_X1 U932 ( .A(n836), .ZN(G319) );
  XOR2_X1 U933 ( .A(G2100), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U934 ( .A(G2090), .B(G2678), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U936 ( .A(n839), .B(KEYINPUT112), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2096), .Z(n843) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1981), .B(G1966), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1961), .B(G1956), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n848), .B(G2474), .Z(n850) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U949 ( .A(KEYINPUT41), .B(G1976), .Z(n852) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1971), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G124), .A2(n875), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n883), .A2(G100), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G136), .A2(n880), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G112), .A2(n876), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n863) );
  XNOR2_X1 U962 ( .A(G164), .B(G160), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n874) );
  NAND2_X1 U964 ( .A1(G106), .A2(n883), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G142), .A2(n880), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT45), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G130), .A2(n875), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G118), .A2(n876), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U971 ( .A(KEYINPUT113), .B(n869), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(G162), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n889) );
  NAND2_X1 U975 ( .A1(G127), .A2(n875), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G115), .A2(n876), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n879), .B(KEYINPUT47), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U981 ( .A1(n883), .A2(G103), .ZN(n884) );
  XOR2_X1 U982 ( .A(KEYINPUT114), .B(n884), .Z(n885) );
  NOR2_X1 U983 ( .A1(n886), .A2(n885), .ZN(n987) );
  XNOR2_X1 U984 ( .A(n887), .B(n987), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U986 ( .A(n972), .B(n890), .Z(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U988 ( .A(n894), .B(n893), .Z(n895) );
  NOR2_X1 U989 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U990 ( .A(n946), .B(KEYINPUT115), .ZN(n897) );
  XNOR2_X1 U991 ( .A(G171), .B(n945), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n900) );
  XNOR2_X1 U993 ( .A(G286), .B(n898), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U995 ( .A1(G37), .A2(n901), .ZN(G397) );
  XNOR2_X1 U996 ( .A(G2451), .B(G2443), .ZN(n911) );
  XOR2_X1 U997 ( .A(G2446), .B(G2454), .Z(n903) );
  XNOR2_X1 U998 ( .A(KEYINPUT110), .B(G2435), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1000 ( .A(KEYINPUT111), .B(G2438), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G2430), .B(G2427), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G57), .ZN(G237) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  XNOR2_X1 U1017 ( .A(G2067), .B(G26), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G32), .B(G1996), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n926) );
  XOR2_X1 U1020 ( .A(G2072), .B(G33), .Z(n921) );
  NAND2_X1 U1021 ( .A1(n921), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G25), .B(n922), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n929) );
  XOR2_X1 U1025 ( .A(G27), .B(n927), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT53), .B(n930), .Z(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(G34), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G2084), .B(n932), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G35), .B(G2090), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n937), .B(KEYINPUT118), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(G29), .A2(n938), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(KEYINPUT55), .B(n939), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(G11), .ZN(n970) );
  XNOR2_X1 U1038 ( .A(G168), .B(G1966), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n941), .B(KEYINPUT120), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(KEYINPUT57), .ZN(n952) );
  XNOR2_X1 U1042 ( .A(n945), .B(G1348), .ZN(n948) );
  XOR2_X1 U1043 ( .A(G1341), .B(n946), .Z(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G1961), .B(G301), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n964) );
  XNOR2_X1 U1048 ( .A(n997), .B(G166), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(KEYINPUT121), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G1956), .B(G299), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(KEYINPUT122), .B(n962), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT119), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT56), .B(n965), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1060 ( .A(KEYINPUT123), .B(n968), .Z(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n996) );
  XOR2_X1 U1062 ( .A(G160), .B(G2084), .Z(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n976) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n981) );
  XOR2_X1 U1066 ( .A(G2090), .B(G162), .Z(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(n979), .B(KEYINPUT51), .ZN(n980) );
  NOR2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1072 ( .A(KEYINPUT116), .B(n986), .ZN(n992) );
  XOR2_X1 U1073 ( .A(G2072), .B(n987), .Z(n989) );
  XOR2_X1 U1074 ( .A(G164), .B(G2078), .Z(n988) );
  NOR2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(KEYINPUT50), .B(n990), .ZN(n991) );
  NAND2_X1 U1077 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(KEYINPUT52), .B(n993), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n994), .A2(G29), .ZN(n995) );
  NAND2_X1 U1080 ( .A1(n996), .A2(n995), .ZN(n1024) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n999) );
  XNOR2_X1 U1082 ( .A(n997), .B(G22), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1085 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(n1002), .Z(n1020) );
  XOR2_X1 U1087 ( .A(G1966), .B(G21), .Z(n1013) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(n1003), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(KEYINPUT125), .B(G1341), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(G19), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  XOR2_X1 U1099 ( .A(KEYINPUT124), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1100 ( .A(G5), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1018), .Z(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1021), .Z(n1022) );
  NOR2_X1 U1105 ( .A1(G16), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1106 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

