//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n468), .B1(new_n461), .B2(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n469), .B2(new_n462), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n465), .B1(new_n470), .B2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n463), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n471), .A2(new_n473), .A3(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT66), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT67), .B1(new_n461), .B2(G2105), .ZN(new_n487));
  AND4_X1   g062(.A1(KEYINPUT67), .A2(new_n471), .A3(new_n473), .A4(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n479), .B1(new_n484), .B2(new_n485), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n471), .A2(new_n473), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n461), .A2(KEYINPUT68), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n462), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n497), .A2(new_n500), .A3(new_n501), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT69), .A3(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(new_n513), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n512), .A2(KEYINPUT69), .A3(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(KEYINPUT69), .B1(new_n512), .B2(G543), .ZN(new_n524));
  OAI211_X1 g099(.A(G62), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(new_n526), .B1(G75), .B2(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n514), .A2(KEYINPUT70), .A3(G62), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n520), .B1(new_n529), .B2(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  AOI211_X1 g106(.A(new_n531), .B(new_n521), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n508), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n526), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT72), .A4(new_n520), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n533), .A2(new_n540), .ZN(G166));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G51), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n519), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n517), .A2(G89), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  AOI22_X1  g125(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n521), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n516), .A2(new_n553), .B1(new_n554), .B2(new_n518), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n511), .A2(new_n513), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(new_n522), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n521), .B1(new_n561), .B2(KEYINPUT74), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(KEYINPUT74), .B2(new_n561), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n517), .A2(G81), .B1(G43), .B2(new_n519), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n519), .A2(G53), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n514), .A2(G91), .A3(new_n515), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n518), .A2(new_n580), .B1(KEYINPUT76), .B2(new_n575), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n514), .A2(G65), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n521), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n582), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  AND2_X1   g162(.A1(new_n533), .A2(new_n540), .ZN(G303));
  NAND4_X1  g163(.A1(new_n558), .A2(G87), .A3(new_n522), .A4(new_n515), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n515), .A2(G49), .A3(G543), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(new_n514), .A2(G61), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n521), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n558), .A2(G86), .A3(new_n522), .A4(new_n515), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n515), .A2(G48), .A3(G543), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n521), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n516), .A2(new_n604), .B1(new_n605), .B2(new_n518), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(G301), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n517), .A2(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n559), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n519), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n618), .A2(KEYINPUT78), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(KEYINPUT78), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n610), .B1(new_n622), .B2(new_n609), .ZN(G284));
  AOI21_X1  g198(.A(new_n610), .B1(new_n622), .B2(new_n609), .ZN(G321));
  NAND2_X1  g199(.A1(G299), .A2(new_n609), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n609), .B2(G168), .ZN(G280));
  XOR2_X1   g201(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g208(.A(new_n484), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G135), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT82), .Z(new_n636));
  INV_X1    g211(.A(new_n489), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n462), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n636), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n482), .A2(G2104), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT81), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n649), .ZN(G156));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n657), .B2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n654), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(G14), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  AOI21_X1  g247(.A(KEYINPUT18), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT85), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n680), .A2(new_n682), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n685), .A3(new_n683), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n688), .B(new_n690), .C1(new_n685), .C2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT33), .ZN(new_n702));
  INV_X1    g277(.A(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G6), .A2(G16), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n600), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G22), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G166), .B2(G16), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n637), .A2(G119), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT87), .B1(G95), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n634), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n718), .B1(new_n727), .B2(new_n717), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n698), .A2(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n607), .B2(new_n698), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1986), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n714), .B2(KEYINPUT34), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G4), .A2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n622), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT88), .B(G1348), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  INV_X1    g319(.A(G139), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n484), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT92), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(new_n462), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2072), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n698), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n566), .B2(new_n698), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT89), .B(G1341), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n742), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n717), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2084), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n698), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n698), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n764), .B1(new_n767), .B2(G1961), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT97), .B(G28), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G168), .A2(new_n698), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n698), .B2(G21), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G2084), .B2(new_n763), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n767), .A2(G1961), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G105), .B2(new_n459), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n634), .A2(G141), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n637), .A2(G129), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n717), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n717), .B2(G32), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT27), .B(G1996), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n780), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G164), .A2(new_n717), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G27), .B2(new_n717), .ZN(new_n795));
  INV_X1    g370(.A(G2078), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n797), .B(new_n798), .C1(new_n641), .C2(new_n717), .ZN(new_n799));
  OR4_X1    g374(.A1(new_n768), .A2(new_n779), .A3(new_n793), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n791), .A2(new_n792), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT95), .ZN(new_n802));
  NAND2_X1  g377(.A1(G299), .A2(G16), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n698), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT23), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G1956), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n776), .A2(new_n777), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  NAND3_X1  g385(.A1(new_n802), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n717), .A2(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G162), .B2(new_n717), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT29), .Z(new_n814));
  INV_X1    g389(.A(G2090), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n717), .A2(G26), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT28), .ZN(new_n818));
  OR2_X1    g393(.A1(G104), .A2(G2105), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n819), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n820));
  INV_X1    g395(.A(G128), .ZN(new_n821));
  INV_X1    g396(.A(G140), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n820), .B1(new_n489), .B2(new_n821), .C1(new_n484), .C2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(new_n717), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT91), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT90), .B(G2067), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n814), .A2(new_n815), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n816), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n758), .A2(new_n800), .A3(new_n811), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n738), .A2(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  AOI22_X1  g408(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n521), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n516), .A2(new_n836), .B1(new_n837), .B2(new_n518), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n839), .A2(new_n842), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n566), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n565), .A2(new_n842), .A3(new_n839), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n622), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT99), .ZN(new_n853));
  INV_X1    g428(.A(G860), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n851), .B2(KEYINPUT39), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n841), .B1(new_n853), .B2(new_n855), .ZN(G145));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n857));
  XNOR2_X1  g432(.A(G160), .B(KEYINPUT100), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT68), .B1(new_n461), .B2(new_n492), .ZN(new_n860));
  AND4_X1   g435(.A1(KEYINPUT68), .A2(new_n471), .A3(new_n473), .A4(new_n492), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n505), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n500), .A2(new_n501), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT101), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n823), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n751), .A2(new_n788), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n634), .A2(G142), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n637), .A2(G130), .ZN(new_n872));
  OR2_X1    g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n789), .A2(new_n748), .A3(new_n750), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n870), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n875), .B1(new_n870), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n869), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n726), .B(new_n646), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n870), .A2(new_n876), .ZN(new_n882));
  INV_X1    g457(.A(new_n875), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n868), .A3(new_n877), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n881), .B1(new_n880), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n859), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n641), .B(G162), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n880), .A2(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(new_n881), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(KEYINPUT102), .A3(new_n886), .A4(new_n858), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n890), .B1(new_n889), .B2(new_n894), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n857), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n894), .ZN(new_n900));
  INV_X1    g475(.A(new_n890), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n896), .A4(new_n895), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n899), .A2(new_n903), .ZN(G395));
  NAND2_X1  g479(.A1(new_n839), .A2(new_n609), .ZN(new_n905));
  NOR2_X1   g480(.A1(G303), .A2(G305), .ZN(new_n906));
  NOR2_X1   g481(.A1(G166), .A2(new_n600), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n607), .B(G288), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT103), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n909), .A2(KEYINPUT103), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n906), .A2(new_n912), .A3(new_n907), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n630), .B(new_n847), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n618), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n618), .A2(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n915), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n905), .B1(new_n927), .B2(new_n609), .ZN(G295));
  OAI21_X1  g503(.A(new_n905), .B1(new_n927), .B2(new_n609), .ZN(G331));
  OR2_X1    g504(.A1(new_n908), .A2(new_n910), .ZN(new_n930));
  INV_X1    g505(.A(new_n913), .ZN(new_n931));
  XNOR2_X1  g506(.A(G286), .B(G171), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n845), .A2(new_n846), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n845), .B2(new_n846), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n922), .B(new_n923), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(new_n918), .A3(new_n917), .A4(new_n933), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n930), .A2(new_n931), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT104), .B1(new_n939), .B2(G37), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n936), .A2(new_n938), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n941), .B(new_n896), .C1(new_n942), .C2(new_n914), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n914), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n939), .A2(G37), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n945), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n944), .B2(new_n945), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g530(.A(KEYINPUT63), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n533), .A2(G8), .A3(new_n540), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n533), .A2(KEYINPUT55), .A3(new_n540), .A4(G8), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n867), .A2(new_n962), .A3(G1384), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n862), .B2(new_n863), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n962), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n482), .A2(G137), .B1(G101), .B2(new_n459), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT65), .B1(new_n475), .B2(G2105), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n466), .B(new_n462), .C1(new_n474), .C2(new_n467), .ZN(new_n969));
  OAI211_X1 g544(.A(G40), .B(new_n967), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n712), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n504), .B1(new_n495), .B2(new_n496), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT101), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT101), .B1(new_n500), .B2(new_n501), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n964), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT107), .B(new_n978), .C1(new_n506), .C2(new_n964), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n971), .B(new_n979), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT108), .B(G2090), .Z(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n973), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT109), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n973), .B(new_n988), .C1(new_n983), .C2(new_n985), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n961), .A2(new_n987), .A3(G8), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT50), .B1(new_n867), .B2(G1384), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n500), .A2(new_n501), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n992), .B2(new_n974), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n970), .B1(new_n978), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n994), .A3(new_n984), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n973), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n959), .B(new_n960), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n977), .A2(G40), .A3(new_n964), .A4(G160), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n592), .A2(G1976), .A3(new_n589), .A4(new_n590), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n591), .A2(new_n1002), .A3(G1976), .A4(new_n592), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(G8), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(G61), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n595), .B1(new_n559), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G651), .ZN(new_n1011));
  INV_X1    g586(.A(new_n599), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n596), .A2(new_n599), .A3(G1981), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n596), .B2(new_n599), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(KEYINPUT49), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(G8), .A3(new_n999), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n703), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n999), .A2(new_n1020), .A3(new_n1004), .A4(G8), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1006), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1006), .A2(new_n1019), .A3(KEYINPUT111), .A4(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n977), .B2(new_n964), .ZN(new_n1027));
  OAI211_X1 g602(.A(G40), .B(G160), .C1(new_n965), .C2(new_n962), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n777), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(G2084), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n983), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G286), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n990), .A2(new_n998), .A3(new_n1026), .A4(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1006), .A2(new_n1021), .A3(new_n1019), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT107), .B1(new_n993), .B2(new_n978), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n965), .A2(new_n981), .A3(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(new_n971), .A3(new_n979), .A4(new_n1030), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n997), .B1(new_n1040), .B2(new_n1029), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1036), .A2(KEYINPUT63), .A3(new_n1041), .A4(G168), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n989), .A2(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n865), .A2(new_n866), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1384), .B1(new_n1044), .B2(new_n974), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n970), .B1(new_n1045), .B2(new_n978), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n1039), .A3(new_n984), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n988), .B1(new_n1047), .B2(new_n973), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1042), .B1(new_n1049), .B2(new_n961), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n959), .B(new_n960), .C1(new_n1043), .C2(new_n1048), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n956), .A2(new_n1035), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1019), .A2(new_n703), .A3(new_n700), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1016), .ZN(new_n1054));
  INV_X1    g629(.A(new_n999), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n997), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n990), .B2(new_n1022), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1035), .A2(new_n956), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1058), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G286), .A2(G8), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT51), .B1(new_n1068), .B2(KEYINPUT120), .ZN(new_n1069));
  OAI211_X1 g644(.A(G8), .B(new_n1069), .C1(new_n1032), .C2(G286), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1068), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1032), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1041), .A2(new_n1071), .A3(new_n1069), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1069), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1033), .A2(new_n1068), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(KEYINPUT121), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n990), .A2(new_n998), .A3(new_n1026), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT122), .B(G1961), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1046), .B2(new_n1039), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n977), .A2(new_n964), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n962), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n970), .B1(KEYINPUT45), .B2(new_n993), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(G2078), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1082), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1083), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n983), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT123), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n977), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n971), .A3(new_n966), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1088), .B1(new_n1098), .B2(G2078), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1080), .A2(new_n1081), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n582), .B2(new_n585), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1097), .A2(new_n971), .A3(new_n966), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1956), .B1(new_n991), .B2(new_n994), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n999), .A2(G2067), .ZN(new_n1112));
  INV_X1    g687(.A(G1348), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n983), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1111), .B1(new_n621), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1105), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1104), .B(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n971), .B1(KEYINPUT50), .B2(new_n965), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n978), .B1(new_n977), .B2(new_n964), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n807), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(new_n1108), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT116), .Z(new_n1123));
  NAND3_X1  g698(.A1(new_n1111), .A2(new_n1121), .A3(KEYINPUT61), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1111), .A2(new_n1121), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT118), .B(KEYINPUT61), .C1(new_n1111), .C2(new_n1121), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1996), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1097), .A2(new_n1131), .A3(new_n971), .A4(new_n966), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n999), .A2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n566), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT61), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(new_n1125), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1138), .B(KEYINPUT59), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1124), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n622), .A2(KEYINPUT60), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(new_n1114), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(KEYINPUT60), .B2(new_n622), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1123), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1093), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT45), .B1(new_n1085), .B2(KEYINPUT105), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(KEYINPUT105), .B2(new_n1085), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n469), .A2(new_n462), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n967), .A2(G40), .A3(new_n1089), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n963), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n983), .A2(KEYINPUT124), .A3(new_n1092), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1154), .A2(new_n1160), .A3(new_n1099), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1152), .B1(new_n1100), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1079), .A2(new_n1164), .A3(new_n1081), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1084), .A2(new_n1090), .A3(new_n1082), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT123), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1167));
  OAI211_X1 g742(.A(G301), .B(new_n1099), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1096), .A2(KEYINPUT125), .A3(G301), .A4(new_n1099), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1152), .B1(new_n1162), .B2(G171), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1165), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1066), .B(new_n1102), .C1(new_n1151), .C2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1156), .A2(new_n970), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n823), .B(G2067), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT106), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n788), .B(new_n1131), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n727), .A2(new_n729), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n727), .A2(new_n729), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n607), .B(G1986), .Z(new_n1186));
  OAI21_X1  g761(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1178), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1189), .A2(new_n1184), .B1(G2067), .B2(new_n823), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1179), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1179), .ZN(new_n1192));
  OR3_X1    g767(.A1(new_n1192), .A2(G1986), .A3(G290), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(KEYINPUT48), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1185), .A2(new_n1179), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT48), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(new_n1193), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1191), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1179), .A2(KEYINPUT46), .A3(new_n1131), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT46), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1192), .B2(G1996), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1181), .A2(new_n789), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1200), .B(new_n1202), .C1(new_n1203), .C2(new_n1192), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT127), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1205), .A2(KEYINPUT47), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(KEYINPUT47), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1199), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1188), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g784(.A1(new_n902), .A2(new_n896), .A3(new_n895), .ZN(new_n1211));
  INV_X1    g785(.A(G319), .ZN(new_n1212));
  NOR4_X1   g786(.A1(G229), .A2(new_n1212), .A3(G401), .A4(G227), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g788(.A1(new_n1214), .A2(new_n954), .ZN(G308));
  OAI211_X1 g789(.A(new_n1211), .B(new_n1213), .C1(new_n952), .C2(new_n953), .ZN(G225));
endmodule


