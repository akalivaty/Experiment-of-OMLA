//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G140), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT80), .B(G110), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT81), .A2(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT81), .A2(G107), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n196), .A2(new_n197), .A3(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT82), .A3(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n198), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n206), .B(G104), .C1(new_n196), .C2(new_n197), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  AND4_X1   g031(.A1(new_n213), .A2(new_n215), .A3(new_n217), .A4(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n216), .B2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT83), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(KEYINPUT1), .C1(new_n216), .C2(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(G128), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n217), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT84), .B1(new_n212), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(G128), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n221), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n218), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n211), .A4(new_n205), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT85), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n242), .A3(G101), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n224), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  INV_X1    g062(.A(new_n224), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n249), .A2(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n253), .B2(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n244), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT10), .B1(new_n226), .B2(new_n233), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT85), .ZN(new_n259));
  INV_X1    g073(.A(new_n212), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n219), .A2(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n224), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n230), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n238), .A2(new_n257), .A3(new_n259), .A4(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n268), .A2(new_n271), .A3(new_n274), .A4(new_n269), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n195), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n264), .B1(new_n258), .B2(KEYINPUT85), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n237), .B(KEYINPUT10), .C1(new_n226), .C2(new_n233), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n276), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(KEYINPUT86), .A3(new_n281), .A4(new_n257), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n265), .A2(new_n276), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n194), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n212), .A2(new_n262), .A3(new_n230), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n234), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(KEYINPUT12), .A3(new_n276), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT12), .B1(new_n287), .B2(new_n276), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n193), .B(new_n290), .C1(new_n277), .C2(new_n282), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n187), .B(new_n188), .C1(new_n285), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n290), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n278), .A2(new_n256), .A3(new_n279), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT86), .B1(new_n294), .B2(new_n281), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n265), .A2(new_n195), .A3(new_n276), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n193), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n193), .B1(new_n277), .B2(new_n282), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n284), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(G469), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(G469), .A2(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n292), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT87), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT2), .B(G113), .ZN(new_n308));
  AND2_X1   g122(.A1(KEYINPUT67), .A2(G116), .ZN(new_n309));
  NOR2_X1   g123(.A1(KEYINPUT67), .A2(G116), .ZN(new_n310));
  OAI21_X1  g124(.A(G119), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT66), .A2(G119), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n308), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT66), .B(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G116), .ZN(new_n321));
  INV_X1    g135(.A(new_n308), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n311), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n241), .A2(new_n324), .A3(new_n243), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT88), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(new_n327), .A3(G116), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n328), .A2(KEYINPUT89), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(KEYINPUT89), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G113), .A3(new_n330), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n312), .A2(new_n318), .A3(new_n327), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n323), .B(new_n260), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n241), .A2(new_n334), .A3(new_n324), .A4(new_n243), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n326), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(G110), .B(G122), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n307), .B1(new_n338), .B2(KEYINPUT6), .ZN(new_n339));
  INV_X1    g153(.A(new_n337), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n326), .A2(new_n340), .A3(new_n333), .A4(new_n335), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(G125), .B2(new_n263), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n189), .A2(G224), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n348), .B(KEYINPUT91), .Z(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n338), .A2(new_n307), .A3(KEYINPUT6), .A4(new_n341), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n331), .B(KEYINPUT92), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n323), .B1(new_n353), .B2(new_n332), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n260), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n323), .B(new_n212), .C1(new_n331), .C2(new_n332), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n337), .B(KEYINPUT8), .Z(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n346), .A2(KEYINPUT93), .B1(KEYINPUT7), .B2(new_n348), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n347), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n359), .A2(new_n347), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n358), .A2(new_n360), .A3(new_n341), .A4(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n352), .A2(new_n188), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G210), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n352), .A2(new_n188), .A3(new_n362), .A4(new_n364), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n306), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT9), .B(G234), .Z(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G221), .B1(new_n370), .B2(G902), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n371), .B(KEYINPUT79), .Z(new_n372));
  XNOR2_X1  g186(.A(G125), .B(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n345), .A2(KEYINPUT16), .A3(G140), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(G146), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT74), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT74), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G146), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n379), .A2(G146), .ZN(new_n383));
  NOR2_X1   g197(.A1(G237), .A2(G953), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(G143), .A3(G214), .ZN(new_n385));
  AOI21_X1  g199(.A(G143), .B1(new_n384), .B2(G214), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT17), .B(G131), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(KEYINPUT95), .A3(new_n383), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n385), .A2(new_n386), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n274), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n390), .A2(KEYINPUT17), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n378), .A2(new_n383), .A3(new_n381), .A4(new_n387), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n200), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n389), .B(new_n398), .Z(new_n399));
  AOI21_X1  g213(.A(KEYINPUT94), .B1(new_n373), .B2(new_n214), .ZN(new_n400));
  OR3_X1    g214(.A1(new_n400), .A2(new_n214), .A3(new_n373), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n214), .B2(new_n373), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n377), .B(KEYINPUT76), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n373), .B(KEYINPUT19), .Z(new_n406));
  OAI211_X1 g220(.A(new_n405), .B(new_n390), .C1(G146), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(new_n397), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G475), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n188), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n395), .A2(new_n397), .A3(new_n403), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n397), .B1(new_n395), .B2(new_n403), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n188), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G475), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n411), .A2(KEYINPUT20), .A3(new_n412), .A4(new_n188), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n422));
  INV_X1    g236(.A(G128), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(G143), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n216), .A2(KEYINPUT96), .A3(G128), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n216), .A2(G128), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n267), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G122), .B1(new_n309), .B2(new_n310), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n196), .A2(new_n197), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g249(.A(KEYINPUT13), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT97), .B1(new_n437), .B2(new_n428), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT13), .B1(new_n424), .B2(new_n425), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(new_n427), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n426), .A2(new_n436), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n429), .B(new_n435), .C1(new_n443), .C2(new_n267), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT98), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n430), .A2(KEYINPUT98), .A3(KEYINPUT14), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n432), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G107), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n430), .A3(new_n432), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n426), .A2(new_n428), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G134), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n429), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G217), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n370), .A2(new_n458), .A3(G953), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n444), .A2(new_n456), .A3(new_n459), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n188), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n464), .B(new_n466), .Z(new_n467));
  NAND2_X1  g281(.A1(new_n421), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G952), .A3(new_n189), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT21), .B(G898), .Z(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n303), .A2(new_n368), .A3(new_n372), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n423), .B1(new_n316), .B2(new_n317), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n315), .A2(G128), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT23), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G110), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n320), .B2(G128), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT75), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT72), .B1(new_n479), .B2(new_n480), .ZN(new_n487));
  INV_X1    g301(.A(new_n317), .ZN(new_n488));
  NOR2_X1   g302(.A1(KEYINPUT66), .A2(G119), .ZN(new_n489));
  OAI21_X1  g303(.A(G128), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n481), .A2(new_n496), .A3(new_n482), .A4(new_n484), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n486), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n373), .A2(new_n214), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n405), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n493), .A2(new_n494), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n378), .A2(new_n383), .A3(new_n381), .ZN(new_n502));
  INV_X1    g316(.A(new_n484), .ZN(new_n503));
  INV_X1    g317(.A(new_n480), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n483), .B1(new_n490), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT73), .B(G110), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n481), .A2(new_n484), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT73), .B1(new_n508), .B2(G110), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n501), .B(new_n502), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n500), .A2(new_n510), .A3(new_n514), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n188), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT77), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT25), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n458), .B1(G234), .B2(new_n188), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT25), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n516), .ZN(new_n526));
  INV_X1    g340(.A(new_n517), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n526), .A2(KEYINPUT78), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n516), .B2(new_n517), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n525), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT64), .ZN(new_n533));
  XNOR2_X1  g347(.A(G134), .B(G137), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n274), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n270), .A2(G134), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n267), .A2(G137), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT64), .B(G131), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n275), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n535), .A2(KEYINPUT69), .A3(new_n538), .A4(new_n275), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n263), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n252), .A2(new_n254), .A3(new_n276), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n312), .A2(new_n318), .A3(new_n308), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n322), .B1(new_n321), .B2(new_n311), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT70), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n324), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT65), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n535), .A2(KEYINPUT65), .A3(new_n538), .A4(new_n275), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n263), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n344), .A2(new_n276), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT28), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n545), .A2(new_n552), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n384), .A2(G210), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n208), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n565), .B(new_n566), .Z(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n567), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n545), .A2(KEYINPUT30), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n557), .A2(new_n571), .A3(new_n558), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n548), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n569), .B1(new_n573), .B2(new_n553), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n545), .A2(new_n552), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n553), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n563), .B1(new_n580), .B2(new_n562), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n567), .A2(KEYINPUT29), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n568), .A2(new_n574), .A3(KEYINPUT71), .A4(new_n575), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n578), .A2(new_n188), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G472), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n557), .A2(new_n571), .A3(new_n558), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n571), .B1(new_n543), .B2(new_n544), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n324), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n561), .A3(new_n567), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n589), .A2(KEYINPUT31), .A3(new_n561), .A4(new_n567), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n560), .A2(new_n563), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n569), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  NOR2_X1   g412(.A1(G472), .A2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n592), .A2(new_n593), .B1(new_n595), .B2(new_n569), .ZN(new_n601));
  INV_X1    g415(.A(new_n599), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT32), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n532), .B1(new_n586), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n478), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n208), .ZN(G3));
  INV_X1    g422(.A(new_n532), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n601), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n597), .A2(new_n599), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n303), .A2(new_n609), .A3(new_n372), .A4(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n372), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n297), .A2(new_n193), .B1(new_n299), .B2(new_n284), .ZN(new_n618));
  OAI21_X1  g432(.A(G469), .B1(new_n618), .B2(G902), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n292), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(KEYINPUT99), .A3(new_n609), .A4(new_n613), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n304), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n366), .B2(new_n367), .ZN(new_n624));
  INV_X1    g438(.A(new_n476), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n464), .A2(new_n465), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n462), .A2(KEYINPUT100), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n444), .A2(new_n456), .A3(new_n629), .A4(new_n459), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n628), .A2(new_n461), .A3(KEYINPUT33), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n630), .A2(KEYINPUT33), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(KEYINPUT101), .A3(new_n461), .A4(new_n628), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n633), .A2(new_n635), .B1(new_n636), .B2(new_n463), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n465), .A2(G902), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n627), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT102), .B1(new_n639), .B2(new_n421), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n635), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n463), .A2(new_n636), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(new_n638), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n626), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n624), .A2(new_n625), .A3(new_n640), .A4(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n622), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NOR2_X1   g466(.A1(new_n467), .A2(new_n646), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n624), .A2(new_n625), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n622), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  AND3_X1   g472(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT25), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n520), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n661), .B(new_n662), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n511), .B(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n660), .A2(new_n522), .B1(new_n525), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n478), .A2(new_n612), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AOI21_X1  g482(.A(new_n665), .B1(new_n586), .B2(new_n604), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n474), .A2(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n470), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n467), .A2(new_n646), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n620), .A2(new_n624), .A3(new_n669), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NAND2_X1  g489(.A1(new_n664), .A2(new_n525), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n524), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n580), .A2(new_n567), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n573), .A2(new_n553), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n567), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n680), .B2(G902), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n677), .B1(new_n604), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT38), .B1(new_n366), .B2(new_n367), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n366), .A2(KEYINPUT38), .A3(new_n367), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n464), .B(new_n466), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n646), .A2(new_n304), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n671), .B(KEYINPUT39), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n620), .A2(KEYINPUT40), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT40), .B1(new_n620), .B2(new_n690), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n682), .B(new_n689), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NOR3_X1   g508(.A1(new_n639), .A2(new_n421), .A3(new_n672), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n620), .A2(new_n624), .A3(new_n669), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OAI21_X1  g511(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n698), .A2(new_n193), .B1(new_n299), .B2(new_n293), .ZN(new_n699));
  OAI21_X1  g513(.A(G469), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n605), .A2(new_n292), .A3(new_n371), .A4(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n648), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT41), .B(G113), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  AND3_X1   g518(.A1(new_n700), .A2(new_n292), .A3(new_n371), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n655), .A2(new_n705), .A3(KEYINPUT105), .A4(new_n605), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n701), .B2(new_n654), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n477), .A3(new_n624), .A4(new_n669), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND3_X1  g526(.A1(new_n700), .A2(new_n292), .A3(new_n371), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n610), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(KEYINPUT106), .B(G472), .C1(new_n601), .C2(G902), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n581), .A2(new_n569), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n602), .B1(new_n594), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n609), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n366), .A2(new_n367), .ZN(new_n722));
  INV_X1    g536(.A(new_n688), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n625), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n713), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n431), .ZN(G24));
  NAND4_X1  g540(.A1(new_n624), .A2(new_n700), .A3(new_n292), .A4(new_n371), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n677), .A3(new_n695), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n345), .ZN(G27));
  AND3_X1   g545(.A1(new_n366), .A2(new_n367), .A3(new_n304), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n303), .A2(new_n732), .A3(new_n371), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n605), .A4(new_n695), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n605), .A2(new_n303), .A3(new_n732), .A4(new_n371), .ZN(new_n736));
  INV_X1    g550(.A(new_n695), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  NAND3_X1  g554(.A1(new_n733), .A2(new_n605), .A3(new_n673), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n743));
  OAI22_X1  g557(.A1(new_n639), .A2(new_n646), .B1(KEYINPUT108), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n745), .B1(new_n644), .B2(new_n421), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n612), .A3(new_n677), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT109), .Z(new_n753));
  AOI21_X1  g567(.A(KEYINPUT45), .B1(new_n298), .B2(new_n300), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT107), .B1(new_n754), .B2(new_n187), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n618), .A2(KEYINPUT45), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(G469), .C1(new_n618), .C2(KEYINPUT45), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n302), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT46), .B1(new_n759), .B2(new_n302), .ZN(new_n761));
  INV_X1    g575(.A(new_n292), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n371), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n732), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n750), .B2(new_n751), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n753), .A2(new_n765), .A3(new_n690), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n763), .B2(new_n764), .ZN(new_n771));
  INV_X1    g585(.A(new_n761), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n302), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n292), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT47), .A3(new_n371), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n586), .A2(new_n604), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n737), .A2(new_n766), .A3(new_n609), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n303), .A2(new_n372), .A3(new_n624), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n669), .A2(new_n673), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n730), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n764), .B1(new_n619), .B2(new_n292), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n688), .B1(new_n366), .B2(new_n367), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n671), .A3(new_n682), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n696), .A4(new_n790), .ZN(new_n791));
  AOI221_X4 g605(.A(new_n719), .B1(new_n524), .B2(new_n676), .C1(new_n715), .C2(new_n716), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n705), .A2(new_n624), .A3(new_n695), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n674), .A3(new_n696), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n788), .A2(new_n792), .A3(new_n695), .A4(new_n732), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n303), .A2(new_n669), .A3(new_n372), .A4(new_n671), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n766), .A2(new_n468), .ZN(new_n802));
  AOI22_X1  g616(.A1(KEYINPUT111), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n800), .A2(KEYINPUT111), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n739), .A2(new_n803), .A3(new_n804), .A4(new_n741), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n666), .A2(new_n607), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n722), .A2(new_n305), .A3(new_n625), .A4(new_n653), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n616), .A2(new_n621), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n639), .A2(new_n421), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n368), .A2(new_n625), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n616), .A2(new_n621), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n702), .A2(new_n725), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n709), .A2(new_n818), .A3(new_n711), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n806), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT53), .B1(new_n799), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n791), .A2(new_n795), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n797), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n805), .A2(new_n816), .A3(new_n819), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n782), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n797), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n796), .B1(new_n791), .B2(new_n795), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n827), .B(KEYINPUT53), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n826), .B1(new_n799), .B2(new_n821), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n825), .A2(new_n835), .A3(KEYINPUT53), .A4(new_n827), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n829), .B1(new_n837), .B2(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n700), .A2(new_n623), .A3(new_n292), .A4(new_n371), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n470), .B1(new_n746), .B2(new_n748), .ZN(new_n843));
  INV_X1    g657(.A(new_n721), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n686), .B1(new_n840), .B2(new_n841), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n366), .A2(KEYINPUT38), .A3(new_n367), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n683), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n623), .A2(new_n700), .A3(new_n292), .A4(new_n371), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(KEYINPUT115), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n747), .B1(new_n744), .B2(new_n745), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n721), .A3(new_n470), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(KEYINPUT50), .A3(new_n853), .A4(new_n842), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n766), .A2(new_n713), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n843), .A3(new_n792), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n604), .A2(new_n681), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n470), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n705), .A2(new_n609), .A3(new_n732), .A4(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n646), .A3(new_n644), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(KEYINPUT116), .A2(new_n855), .A3(new_n857), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n847), .B2(new_n854), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT116), .B1(new_n864), .B2(new_n857), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n700), .A2(new_n292), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n617), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n771), .A2(new_n775), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n732), .A3(new_n853), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT117), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n864), .A2(new_n857), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(KEYINPUT51), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n856), .A2(new_n843), .A3(new_n605), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT48), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n640), .A2(new_n647), .ZN(new_n878));
  OAI211_X1 g692(.A(G952), .B(new_n189), .C1(new_n860), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n853), .A2(new_n624), .A3(new_n705), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n871), .A2(KEYINPUT117), .A3(new_n872), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n838), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(G952), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n189), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n867), .B(KEYINPUT49), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n849), .A2(new_n617), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n858), .A2(new_n532), .A3(new_n646), .A4(new_n639), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n889), .A2(new_n305), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n892), .ZN(G75));
  NAND2_X1  g707(.A1(new_n886), .A2(G953), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT118), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n822), .A2(new_n828), .A3(G902), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n343), .A2(new_n351), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n350), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n903), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n896), .B1(new_n904), .B2(new_n906), .ZN(G51));
  AND3_X1   g721(.A1(new_n822), .A2(new_n828), .A3(new_n782), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(new_n829), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n302), .B(KEYINPUT57), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n909), .A2(new_n910), .B1(new_n285), .B2(new_n291), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n759), .B(KEYINPUT119), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n897), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n896), .B1(new_n911), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(new_n411), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n411), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n896), .B1(new_n916), .B2(new_n917), .ZN(G60));
  INV_X1    g732(.A(new_n637), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n838), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n921), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n637), .B(new_n923), .C1(new_n908), .C2(new_n829), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n922), .A2(new_n895), .A3(new_n924), .ZN(G63));
  AND2_X1   g739(.A1(new_n822), .A2(new_n828), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n528), .A2(new_n530), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n664), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n895), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n895), .A3(new_n932), .A4(new_n934), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(G66));
  NAND2_X1  g752(.A1(new_n817), .A2(new_n820), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n189), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT121), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n189), .B1(new_n472), .B2(G224), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n901), .B1(G898), .B2(new_n189), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT122), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  AND2_X1   g760(.A1(new_n786), .A2(new_n696), .ZN(new_n947));
  NAND2_X1  g761(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n947), .A2(new_n693), .A3(new_n948), .ZN(new_n949));
  OR2_X1    g763(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n950));
  AOI22_X1  g764(.A1(new_n947), .A2(new_n693), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n813), .A2(new_n653), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n606), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(new_n620), .A3(new_n690), .A4(new_n732), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n780), .A2(new_n952), .A3(new_n768), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n189), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n570), .A2(new_n572), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n406), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(G900), .B2(G953), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n765), .A2(new_n605), .A3(new_n690), .A4(new_n789), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n947), .A2(new_n739), .A3(new_n741), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n780), .A2(new_n768), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(G953), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n966), .B(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n956), .B2(new_n939), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n679), .B(KEYINPUT126), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n569), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n973), .A2(KEYINPUT127), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT127), .B1(new_n973), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n972), .B1(new_n964), .B2(new_n939), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n569), .A3(new_n974), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n895), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n574), .A2(new_n590), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n837), .A2(new_n972), .A3(new_n982), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(G57));
endmodule


