//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT66), .B(G244), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n207), .A2(G77), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G107), .A2(G264), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n206), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n215), .B(new_n218), .C1(new_n221), .C2(new_n223), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT2), .B(G226), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n228), .B(new_n231), .Z(G358));
  XNOR2_X1  g0032(.A(G50), .B(G68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(new_n234));
  XOR2_X1   g0034(.A(G58), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G169), .ZN(new_n241));
  OR2_X1    g0041(.A1(G223), .A2(G1698), .ZN(new_n242));
  INV_X1    g0042(.A(G226), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G1698), .ZN(new_n244));
  AND2_X1   g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NOR2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  OAI211_X1 g0046(.A(new_n242), .B(new_n244), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G87), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(new_n251), .A3(G274), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n251), .A2(G232), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n241), .B1(new_n253), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n251), .B1(new_n247), .B2(new_n248), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n260), .ZN(new_n264));
  INV_X1    g0064(.A(G179), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT16), .ZN(new_n268));
  INV_X1    g0068(.A(G68), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n245), .A2(new_n246), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n219), .A3(KEYINPUT7), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n269), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G58), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n269), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G58), .A2(G68), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G159), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n268), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n220), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT78), .B1(new_n245), .B2(new_n246), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT78), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n274), .A2(new_n292), .A3(new_n276), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n291), .A2(new_n293), .A3(new_n278), .A4(new_n219), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n269), .B1(new_n277), .B2(KEYINPUT7), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n287), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(KEYINPUT16), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n288), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n290), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n302), .A2(new_n275), .A3(G1), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n258), .A2(G20), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT71), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT8), .B(G58), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n304), .A2(new_n308), .B1(new_n303), .B2(new_n307), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n267), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT18), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n253), .A2(new_n261), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n263), .B2(new_n264), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n299), .A2(new_n309), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n274), .A2(new_n276), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(G222), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(G223), .A3(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n270), .A2(G77), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT69), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n251), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT69), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n251), .A2(new_n259), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n257), .B1(new_n243), .B2(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(new_n265), .ZN(new_n336));
  INV_X1    g0136(.A(G50), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n306), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n304), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n285), .A2(G150), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n219), .A2(G33), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n340), .B1(new_n275), .B2(new_n201), .C1(new_n341), .C2(new_n307), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n301), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n303), .A2(new_n337), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n328), .A2(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n336), .B(new_n345), .C1(G169), .C2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n302), .A2(G1), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G20), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G77), .ZN(new_n350));
  INV_X1    g0150(.A(new_n290), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT74), .B1(new_n351), .B2(new_n349), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n303), .A2(new_n290), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n306), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n350), .B1(new_n356), .B2(G77), .ZN(new_n357));
  INV_X1    g0157(.A(new_n285), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n202), .A2(new_n219), .B1(new_n307), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n362), .B(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n361), .B1(new_n364), .B2(new_n341), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n359), .A2(new_n360), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n290), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n321), .A2(G232), .A3(new_n322), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n321), .A2(G238), .A3(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G107), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n321), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n252), .ZN(new_n373));
  INV_X1    g0173(.A(new_n331), .ZN(new_n374));
  INV_X1    g0174(.A(G274), .ZN(new_n375));
  AND2_X1   g0175(.A1(G1), .A2(G13), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n250), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n374), .A2(new_n207), .B1(new_n256), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n241), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(new_n265), .A3(new_n378), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n368), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(G200), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n373), .A2(G190), .A3(new_n378), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(new_n357), .A3(new_n367), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n347), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n312), .A2(new_n320), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n330), .A2(new_n335), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT9), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n345), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT9), .A4(new_n344), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n388), .A2(new_n313), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n391), .A2(new_n392), .ZN(new_n396));
  INV_X1    g0196(.A(new_n394), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT10), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n389), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT79), .ZN(new_n402));
  INV_X1    g0202(.A(G238), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n257), .B1(new_n403), .B2(new_n331), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n321), .A2(G226), .A3(new_n322), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT75), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT75), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(G33), .A3(G97), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(G232), .B(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(KEYINPUT13), .B(new_n404), .C1(new_n252), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n252), .ZN(new_n415));
  INV_X1    g0215(.A(new_n404), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(G169), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(KEYINPUT76), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT76), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n404), .B1(new_n412), .B2(new_n252), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(new_n414), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n414), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n420), .A2(G179), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(G169), .C1(new_n413), .C2(new_n417), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n356), .A2(G68), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n269), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n341), .B2(new_n202), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n301), .A3(KEYINPUT11), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n301), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT11), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n303), .A2(new_n269), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT12), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n429), .A2(new_n432), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n413), .A2(new_n417), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n440), .B2(G200), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n313), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n443), .A3(KEYINPUT77), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n439), .A2(new_n443), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n401), .A2(new_n402), .A3(new_n444), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n444), .A3(new_n400), .A4(new_n387), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n403), .A2(new_n322), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n453), .B1(G244), .B2(new_n322), .C1(new_n245), .C2(new_n246), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n251), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n251), .A2(G274), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n258), .A2(G45), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G250), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n457), .A2(new_n458), .B1(new_n252), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G179), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n241), .B2(new_n461), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n362), .B(KEYINPUT73), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n349), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n219), .B1(new_n410), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G87), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n371), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n472), .A2(new_n474), .A3(G33), .A4(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n321), .A2(new_n219), .A3(G68), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(new_n479), .A3(new_n466), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n471), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n465), .B1(new_n481), .B2(new_n290), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n290), .B(KEYINPUT70), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT81), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n273), .B2(G1), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n258), .A2(KEYINPUT81), .A3(G33), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n483), .A2(new_n349), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n464), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT85), .B1(new_n482), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n463), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(G200), .B1(new_n456), .B2(new_n460), .ZN(new_n495));
  INV_X1    g0295(.A(new_n460), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n454), .A2(new_n455), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n251), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n313), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(G244), .B(new_n322), .C1(new_n245), .C2(new_n246), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n321), .A2(KEYINPUT4), .A3(G244), .A4(new_n322), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n321), .A2(G250), .A3(G1698), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n252), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n255), .A2(G1), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n254), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(G41), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n377), .A2(new_n510), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n510), .A3(new_n511), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n251), .ZN(new_n517));
  INV_X1    g0317(.A(G257), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n241), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT7), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n371), .B1(new_n202), .B2(new_n358), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT80), .B(G107), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n469), .A2(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n469), .A2(new_n371), .A3(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n529), .A3(new_n528), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n219), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n290), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n349), .A2(G97), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n488), .B2(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n519), .B1(new_n252), .B2(new_n508), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT83), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(new_n265), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n538), .B2(new_n265), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n522), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n472), .B(new_n474), .C1(new_n245), .C2(new_n246), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT22), .B1(new_n543), .B2(new_n468), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n321), .A2(new_n219), .A3(new_n545), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT23), .A2(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(G20), .ZN(new_n551));
  INV_X1    g0351(.A(new_n219), .ZN(new_n552));
  NOR2_X1   g0352(.A1(KEYINPUT23), .A2(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n548), .B1(new_n547), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n290), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n303), .A2(new_n371), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT25), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n488), .B2(G107), .ZN(new_n561));
  OAI211_X1 g0361(.A(G257), .B(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n562));
  OAI211_X1 g0362(.A(G250), .B(new_n322), .C1(new_n245), .C2(new_n246), .ZN(new_n563));
  INV_X1    g0363(.A(G294), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n273), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n252), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n516), .A2(G264), .A3(new_n251), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n515), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G190), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT90), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n516), .A2(KEYINPUT90), .A3(G264), .A4(new_n251), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n252), .B2(new_n565), .ZN(new_n573));
  AOI21_X1  g0373(.A(G200), .B1(new_n573), .B2(new_n515), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n558), .B(new_n561), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n271), .A2(new_n279), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G107), .B1(G77), .B2(new_n285), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n531), .A2(new_n532), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n552), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n351), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n535), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n483), .A2(new_n349), .A3(new_n487), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n469), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n538), .A2(G190), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n521), .A2(G200), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n542), .A2(new_n575), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n547), .A2(new_n554), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n351), .B1(new_n590), .B2(new_n555), .ZN(new_n591));
  INV_X1    g0391(.A(new_n561), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT89), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT89), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n558), .A2(new_n594), .A3(new_n561), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n568), .A2(G169), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n573), .A2(new_n515), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n265), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n516), .A2(G270), .A3(new_n251), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n515), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G257), .B(new_n322), .C1(new_n245), .C2(new_n246), .ZN(new_n603));
  OAI211_X1 g0403(.A(G264), .B(G1698), .C1(new_n245), .C2(new_n246), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n274), .A2(G303), .A3(new_n276), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n252), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(KEYINPUT21), .A3(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n265), .B2(new_n608), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n219), .B(new_n506), .C1(G33), .C2(new_n469), .ZN(new_n611));
  INV_X1    g0411(.A(G116), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n289), .A2(new_n220), .B1(G20), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(KEYINPUT87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(KEYINPUT87), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(G116), .B(new_n487), .C1(new_n352), .C2(new_n354), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n303), .A2(new_n612), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT86), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n611), .A2(KEYINPUT87), .A3(new_n615), .A4(new_n613), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n618), .A2(new_n619), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G169), .A3(new_n608), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n610), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n606), .A2(new_n252), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n627), .A2(G190), .A3(new_n601), .ZN(new_n628));
  AOI21_X1  g0428(.A(G200), .B1(new_n602), .B2(new_n607), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT88), .B1(new_n630), .B2(new_n623), .ZN(new_n631));
  INV_X1    g0431(.A(new_n623), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT88), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(new_n633), .C1(new_n628), .C2(new_n629), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n599), .A2(new_n626), .A3(new_n635), .ZN(new_n636));
  NOR4_X1   g0436(.A1(new_n452), .A2(new_n501), .A3(new_n588), .A4(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n481), .A2(new_n290), .ZN(new_n638));
  INV_X1    g0438(.A(new_n465), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(new_n489), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n463), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n495), .A2(KEYINPUT91), .B1(new_n461), .B2(G190), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n498), .A2(new_n643), .A3(G200), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n642), .A2(new_n482), .A3(new_n493), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT92), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT92), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n580), .A2(new_n583), .B1(G169), .B2(new_n538), .ZN(new_n652));
  INV_X1    g0452(.A(new_n541), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n538), .A2(new_n539), .A3(new_n265), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n542), .A2(new_n575), .A3(new_n587), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n598), .B1(new_n591), .B2(new_n592), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n626), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n650), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n641), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n492), .A2(new_n655), .A3(new_n500), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n656), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n451), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT93), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT93), .B1(new_n395), .B2(new_n399), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n382), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n443), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n439), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n318), .B(KEYINPUT17), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n312), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n347), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n665), .A2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n610), .A2(new_n623), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n625), .A2(new_n624), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n219), .A2(new_n348), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT95), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n593), .A2(new_n595), .A3(new_n687), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n599), .A2(new_n691), .A3(new_n575), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n599), .B2(new_n688), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n658), .A2(new_n687), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n632), .A2(new_n688), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n681), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n635), .A2(new_n626), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(KEYINPUT94), .B(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n693), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(G399));
  NAND2_X1  g0505(.A1(new_n216), .A2(new_n254), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n470), .A2(G116), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n707), .A2(new_n258), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n223), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  NAND2_X1  g0511(.A1(new_n662), .A2(new_n651), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n641), .A2(new_n645), .A3(new_n648), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n648), .B1(new_n641), .B2(new_n645), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT26), .B(new_n655), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n599), .A2(new_n626), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n650), .A2(new_n717), .A3(new_n657), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n641), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .A3(new_n688), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT99), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n588), .B1(new_n649), .B2(new_n647), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n661), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n687), .B1(new_n723), .B2(new_n716), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT99), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT29), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n664), .A2(new_n688), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n721), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n573), .A2(new_n461), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n608), .A2(new_n265), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT97), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n731), .A2(new_n538), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n627), .A2(new_n601), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n538), .A2(new_n737), .A3(G179), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n734), .B1(new_n738), .B2(new_n730), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n737), .A2(G179), .A3(new_n461), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n573), .A2(new_n515), .B1(new_n509), .B2(new_n520), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(KEYINPUT98), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n597), .A2(KEYINPUT98), .A3(new_n521), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n736), .B(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n687), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT96), .B(KEYINPUT31), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n702), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n636), .ZN(new_n749));
  INV_X1    g0549(.A(new_n501), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n657), .A4(new_n688), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n745), .A2(KEYINPUT31), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n729), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n711), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n552), .A2(new_n302), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G45), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G1), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n707), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n703), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n702), .B2(new_n700), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n216), .A2(G355), .A3(new_n321), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G116), .B2(new_n216), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n236), .A2(new_n255), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n291), .A2(new_n293), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n216), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n255), .B2(new_n223), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n220), .B1(G20), .B2(new_n241), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n759), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n275), .A2(new_n313), .A3(new_n315), .A4(G179), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n270), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n219), .A2(new_n265), .A3(G190), .A4(new_n315), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT33), .B(G317), .Z(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n552), .B1(new_n313), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n781), .A2(new_n782), .B1(new_n786), .B2(new_n564), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n219), .A2(new_n265), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G190), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n779), .B(new_n787), .C1(G311), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(G190), .A3(new_n315), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT101), .B(G326), .Z(new_n797));
  AOI22_X1  g0597(.A1(G322), .A2(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n219), .A2(G190), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT100), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n784), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G329), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n800), .A2(G179), .A3(new_n315), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G283), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n792), .A2(new_n798), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(G159), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n803), .A2(G107), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n777), .A2(new_n468), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n270), .B(new_n809), .C1(new_n780), .C2(G68), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n786), .A2(new_n469), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G77), .B2(new_n791), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G50), .A2(new_n796), .B1(new_n794), .B2(G58), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n808), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n805), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n775), .B1(new_n772), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n771), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n700), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n761), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NOR2_X1   g0620(.A1(new_n382), .A2(new_n687), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n368), .A2(new_n687), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n385), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n382), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n728), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n826), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n664), .A2(new_n688), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n753), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(KEYINPUT104), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(KEYINPUT104), .ZN(new_n833));
  INV_X1    g0633(.A(new_n759), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n827), .A2(new_n753), .A3(new_n829), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n828), .A2(new_n770), .ZN(new_n837));
  INV_X1    g0637(.A(new_n772), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n770), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n781), .A2(new_n840), .B1(new_n612), .B2(new_n790), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n841), .A2(KEYINPUT102), .B1(G303), .B2(new_n796), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(KEYINPUT102), .B2(new_n841), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT103), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n803), .A2(G87), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n321), .B(new_n811), .C1(G107), .C2(new_n776), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n801), .A2(G311), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n794), .A2(G294), .ZN(new_n848));
  AND4_X1   g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n791), .A2(G159), .B1(G150), .B2(new_n780), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  INV_X1    g0651(.A(G143), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n851), .B2(new_n795), .C1(new_n852), .C2(new_n793), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT34), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n803), .A2(G68), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n765), .B1(G50), .B2(new_n776), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(new_n281), .C2(new_n786), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G132), .B2(new_n801), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n844), .A2(new_n849), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n759), .B1(G77), .B2(new_n839), .C1(new_n859), .C2(new_n838), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n832), .A2(new_n836), .B1(new_n837), .B2(new_n860), .ZN(G384));
  OAI21_X1  g0661(.A(G77), .B1(new_n281), .B2(new_n269), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n862), .A2(new_n222), .B1(G50), .B2(new_n269), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(G1), .A3(new_n302), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT105), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n221), .A2(G116), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n578), .B2(KEYINPUT35), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(KEYINPUT35), .B2(new_n578), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT36), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n829), .A2(new_n822), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n299), .A2(new_n309), .ZN(new_n873));
  INV_X1    g0673(.A(new_n267), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n685), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(new_n877), .A3(new_n878), .A4(new_n318), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT106), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n299), .A2(new_n309), .A3(new_n317), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n310), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT106), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n878), .A4(new_n877), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n298), .A2(new_n301), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n296), .B2(new_n297), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n309), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n874), .B2(new_n876), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n878), .B1(new_n889), .B2(new_n318), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n876), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n310), .B(KEYINPUT18), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n674), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n890), .B1(new_n880), .B2(new_n884), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n895), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n438), .A2(new_n687), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n439), .A2(new_n443), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n902), .B1(new_n439), .B2(new_n443), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n872), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n894), .A2(new_n876), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n439), .A2(new_n687), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT107), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  AOI211_X1 g0715(.A(KEYINPUT107), .B(new_n915), .C1(new_n897), .C2(new_n900), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n877), .B1(new_n894), .B2(new_n674), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n685), .B1(new_n299), .B2(new_n309), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n881), .A2(new_n310), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n878), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n885), .B2(KEYINPUT108), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT108), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n880), .A2(new_n884), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n917), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n897), .B1(new_n924), .B2(KEYINPUT38), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n914), .A2(new_n916), .B1(new_n925), .B2(KEYINPUT39), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n911), .B1(new_n912), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n721), .A2(new_n726), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n448), .A2(new_n450), .B1(new_n728), .B2(new_n727), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n676), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n927), .B(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n828), .B1(new_n904), .B2(new_n905), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT109), .ZN(new_n934));
  NOR4_X1   g0734(.A1(new_n636), .A2(new_n501), .A3(new_n588), .A4(new_n687), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n936));
  INV_X1    g0736(.A(new_n743), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n741), .A2(KEYINPUT98), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n937), .A2(new_n938), .A3(new_n740), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n736), .A2(new_n739), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n688), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n936), .B1(new_n941), .B2(new_n747), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n934), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n747), .B1(new_n744), .B2(new_n687), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n751), .A2(new_n946), .A3(KEYINPUT109), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n932), .B(new_n933), .C1(new_n943), .C2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n933), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n935), .A2(new_n942), .A3(new_n934), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT109), .B1(new_n751), .B2(new_n946), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n901), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n948), .A2(new_n925), .B1(new_n952), .B2(new_n932), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n451), .B1(new_n951), .B2(new_n950), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n701), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n931), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n258), .B2(new_n756), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n931), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n871), .B1(new_n959), .B2(new_n960), .ZN(G367));
  NOR2_X1   g0761(.A1(new_n766), .A2(new_n231), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n773), .B1(new_n364), .B2(new_n216), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n803), .A2(G97), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n791), .A2(G283), .B1(G294), .B2(new_n780), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n371), .C2(new_n786), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n777), .A2(new_n612), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT46), .ZN(new_n968));
  INV_X1    g0768(.A(new_n765), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n967), .B2(KEYINPUT46), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(G311), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n971), .B1(new_n778), .B2(new_n793), .C1(new_n972), .C2(new_n795), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n966), .B(new_n973), .C1(G317), .C2(new_n801), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n803), .A2(G77), .ZN(new_n975));
  INV_X1    g0775(.A(new_n801), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n851), .B2(new_n976), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n321), .B1(new_n777), .B2(new_n281), .C1(new_n786), .C2(new_n269), .ZN(new_n978));
  INV_X1    g0778(.A(G159), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n781), .A2(new_n979), .B1(new_n337), .B2(new_n790), .ZN(new_n980));
  INV_X1    g0780(.A(G150), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n852), .A2(new_n795), .B1(new_n793), .B2(new_n981), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n977), .A2(new_n978), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n974), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n759), .B1(new_n962), .B2(new_n963), .C1(new_n985), .C2(new_n838), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n494), .A2(new_n687), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n650), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n641), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n986), .B1(new_n771), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT111), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n542), .A2(new_n688), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT110), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n542), .B(new_n587), .C1(new_n584), .C2(new_n688), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT45), .B1(new_n696), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n996), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n694), .A2(new_n998), .A3(new_n999), .A4(new_n695), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n696), .B2(new_n996), .ZN(new_n1003));
  OAI211_X1 g0803(.A(KEYINPUT44), .B(new_n998), .C1(new_n694), .C2(new_n695), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n703), .B(new_n693), .C1(new_n1001), .C2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n704), .C1(new_n1000), .C2(new_n997), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n703), .B(new_n693), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n690), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n754), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n754), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n706), .B(KEYINPUT41), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n758), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n542), .B1(new_n998), .B2(new_n599), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n694), .A2(new_n996), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n688), .A2(new_n1017), .B1(new_n1018), .B2(KEYINPUT42), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(KEYINPUT42), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n990), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(new_n1020), .B1(KEYINPUT43), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n990), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1022), .B(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n704), .A2(new_n998), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1025), .B(new_n1026), .Z(new_n1027));
  OAI21_X1  g0827(.A(new_n992), .B1(new_n1016), .B2(new_n1027), .ZN(G387));
  OR2_X1    g0828(.A1(new_n693), .A2(new_n817), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n791), .A2(G303), .B1(G311), .B2(new_n780), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  INV_X1    g0831(.A(G322), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n793), .C1(new_n1032), .C2(new_n795), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n785), .A2(G283), .B1(new_n776), .B2(G294), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n803), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n612), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n969), .B(new_n1043), .C1(new_n801), .C2(new_n797), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n781), .A2(new_n307), .B1(new_n269), .B2(new_n790), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n969), .B1(new_n202), .B2(new_n777), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n786), .A2(new_n364), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G50), .A2(new_n794), .B1(new_n796), .B2(G159), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n801), .A2(G150), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n964), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n838), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n216), .A2(new_n321), .A3(new_n708), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(G107), .B2(new_n216), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n228), .A2(G45), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT112), .ZN(new_n1057));
  AOI211_X1 g0857(.A(G45), .B(new_n708), .C1(G68), .C2(G77), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n307), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n766), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1055), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n774), .B1(new_n1063), .B2(KEYINPUT113), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n834), .B(new_n1053), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1011), .A2(new_n758), .B1(new_n1029), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1012), .A2(new_n707), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n754), .A2(new_n1011), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  INV_X1    g0870(.A(new_n758), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n996), .A2(new_n817), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT114), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n773), .B1(new_n469), .B2(new_n216), .C1(new_n766), .C2(new_n239), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n981), .A2(new_n795), .B1(new_n793), .B2(new_n979), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT51), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n969), .B1(new_n269), .B2(new_n777), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G50), .B2(new_n780), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n786), .A2(new_n202), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n307), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n791), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n845), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1076), .B(new_n1082), .C1(G143), .C2(new_n801), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n801), .A2(G322), .B1(G283), .B2(new_n776), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT116), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n786), .A2(new_n612), .B1(new_n564), .B2(new_n790), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n321), .B(new_n1086), .C1(G303), .C2(new_n780), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n972), .A2(new_n793), .B1(new_n795), .B2(new_n1031), .ZN(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1087), .A2(new_n808), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1083), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n759), .B(new_n1074), .C1(new_n1094), .C2(new_n838), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1009), .A2(new_n1071), .B1(new_n1073), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n707), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G390));
  NOR2_X1   g0900(.A1(new_n720), .A2(KEYINPUT99), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n725), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n929), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G330), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n943), .B2(new_n947), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n451), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n677), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n930), .A2(new_n1109), .A3(new_n1106), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n907), .B1(new_n753), .B2(new_n828), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n949), .B2(new_n1105), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n872), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n907), .B1(new_n1105), .B2(new_n828), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n821), .B1(new_n724), .B2(new_n825), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n753), .A2(new_n828), .A3(new_n907), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1108), .A2(new_n1110), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n912), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1120), .B(new_n925), .C1(new_n1115), .C2(new_n906), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n912), .B1(new_n872), .B2(new_n907), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1116), .C1(new_n926), .C2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n883), .B1(new_n919), .B2(new_n878), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n879), .A2(KEYINPUT106), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT108), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n920), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n923), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n917), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT38), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n899), .A2(new_n898), .A3(new_n895), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1120), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n719), .A2(new_n688), .A3(new_n825), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n906), .B1(new_n1133), .B2(new_n822), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT38), .B1(new_n892), .B2(new_n896), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT39), .B1(new_n1136), .B2(new_n1131), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT107), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n901), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1131), .B1(new_n1140), .B2(new_n898), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1138), .A2(new_n1139), .B1(new_n1141), .B2(new_n915), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1122), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1105), .A2(new_n949), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1123), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1119), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n706), .B1(new_n1119), .B2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1146), .A2(new_n1071), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n759), .B1(new_n1080), .B2(new_n839), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n781), .A2(new_n371), .B1(new_n469), .B2(new_n790), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1152), .A2(new_n1079), .A3(new_n321), .A4(new_n809), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G116), .A2(new_n794), .B1(new_n796), .B2(G283), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n801), .A2(G294), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1153), .A2(new_n855), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G125), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n321), .B1(new_n976), .B2(new_n1157), .C1(new_n1042), .C2(new_n337), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT118), .Z(new_n1159));
  OR3_X1    g0959(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n981), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT53), .B1(new_n777), .B2(new_n981), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n781), .C2(new_n851), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT54), .B(G143), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n786), .A2(new_n979), .B1(new_n790), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  INV_X1    g0966(.A(G132), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n795), .C1(new_n1167), .C2(new_n793), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1156), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1151), .B1(new_n1169), .B2(new_n772), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n926), .B2(new_n770), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1149), .A2(new_n1150), .A3(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n952), .A2(new_n932), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n933), .B1(new_n943), .B2(new_n947), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n925), .A2(new_n1174), .A3(KEYINPUT40), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1175), .A3(G330), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n345), .A2(new_n876), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n669), .B2(new_n347), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT93), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n400), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n347), .A3(new_n666), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1179), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1178), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n669), .A2(new_n347), .A3(new_n1179), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n1177), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1176), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1173), .A2(new_n1190), .A3(new_n1175), .A4(G330), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n908), .B(new_n910), .C1(new_n1142), .C2(new_n1120), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT124), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1190), .B1(new_n953), .B2(G330), .ZN(new_n1197));
  AND4_X1   g0997(.A1(G330), .A2(new_n1173), .A3(new_n1190), .A4(new_n1175), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1192), .A2(new_n927), .A3(new_n1193), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1196), .B1(new_n1201), .B2(KEYINPUT124), .ZN(new_n1202));
  AND4_X1   g1002(.A1(new_n1109), .A2(new_n1103), .A3(new_n677), .A4(new_n1106), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1109), .B1(new_n930), .B2(new_n1106), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1118), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1146), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT57), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n707), .B1(new_n1202), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1201), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n759), .B1(G50), .B2(new_n839), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n786), .A2(new_n981), .B1(new_n777), .B2(new_n1163), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n781), .A2(new_n1167), .B1(new_n851), .B2(new_n790), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1157), .A2(new_n795), .B1(new_n793), .B2(new_n1166), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n801), .A2(G124), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G33), .A2(G41), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT119), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n803), .B2(G159), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n803), .A2(G58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n801), .A2(G283), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n791), .A2(new_n464), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n765), .A2(new_n254), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G97), .B2(new_n780), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n785), .A2(G68), .B1(new_n776), .B2(G77), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n795), .B2(new_n612), .C1(new_n371), .C2(new_n793), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT120), .Z(new_n1234));
  XNOR2_X1  g1034(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1228), .A2(new_n337), .A3(new_n1222), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1238), .A2(KEYINPUT122), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(KEYINPUT122), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1224), .B1(new_n1234), .B2(new_n1235), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1212), .B1(new_n1241), .B2(new_n772), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n770), .B2(new_n1190), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT123), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1201), .B2(new_n758), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1211), .A2(new_n1245), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n1118), .A2(new_n758), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n759), .B1(G68), .B2(new_n839), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n969), .B1(new_n979), .B2(new_n777), .C1(new_n790), .C2(new_n981), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n781), .A2(new_n1163), .B1(new_n786), .B2(new_n337), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n1167), .B2(new_n795), .C1(new_n851), .C2(new_n793), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1225), .B1(new_n1166), .B2(new_n976), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n321), .B(new_n1048), .C1(G97), .C2(new_n776), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n791), .A2(G107), .B1(G116), .B2(new_n780), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G283), .A2(new_n794), .B1(new_n796), .B2(G294), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n975), .B1(new_n778), .B2(new_n976), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1252), .A2(new_n1253), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1248), .B1(new_n1259), .B2(new_n772), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n907), .B2(new_n770), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1247), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1119), .A2(new_n1015), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1118), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(G381));
  NOR2_X1   g1066(.A1(G375), .A2(G378), .ZN(new_n1267));
  INV_X1    g1067(.A(G390), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1271), .A2(G387), .A3(G381), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1273), .A2(KEYINPUT125), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(KEYINPUT125), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G407));
  INV_X1    g1076(.A(G213), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1267), .B2(new_n686), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1274), .B2(new_n1275), .ZN(G409));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1119), .A2(new_n707), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1265), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1206), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT60), .B1(new_n1286), .B2(KEYINPUT126), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1282), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(G384), .A3(new_n1263), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1284), .B1(new_n1265), .B2(new_n1283), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1286), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1281), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1269), .B1(new_n1292), .B2(new_n1262), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1277), .A2(G343), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G2897), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1289), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G378), .B(new_n1245), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1149), .A2(new_n1150), .A3(new_n1171), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1207), .A2(new_n1015), .A3(new_n1201), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1303), .B(new_n1243), .C1(new_n1202), .C2(new_n1071), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1295), .B1(new_n1301), .B2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1280), .B1(new_n1300), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1295), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1294), .ZN(new_n1311));
  AND4_X1   g1111(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1308), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1307), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G387), .A2(new_n1268), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(G393), .B(new_n819), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G390), .B(new_n992), .C1(new_n1016), .C2(new_n1027), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1316), .B1(new_n1315), .B2(new_n1317), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1289), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1296), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1325), .A2(new_n1320), .A3(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1309), .A2(new_n1311), .A3(KEYINPUT63), .A4(new_n1310), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT127), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1306), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1311), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  OAI22_X1  g1134(.A1(new_n1314), .A2(new_n1320), .B1(new_n1329), .B2(new_n1334), .ZN(G405));
  AOI21_X1  g1135(.A(G378), .B1(new_n1211), .B2(new_n1245), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1301), .ZN(new_n1337));
  OR3_X1    g1137(.A1(new_n1336), .A2(new_n1337), .A3(new_n1311), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1311), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1320), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1338), .A2(new_n1320), .A3(new_n1339), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(G402));
endmodule


