//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  OR3_X1    g0004(.A1(new_n204), .A2(KEYINPUT65), .A3(G13), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT65), .B1(new_n204), .B2(G13), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G107), .C2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n204), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(G58), .A2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n209), .B(new_n230), .C1(new_n233), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(G270), .Z(new_n241));
  XOR2_X1   g0041(.A(G238), .B(G244), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G226), .B(G232), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n241), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n264), .B(new_n266), .C1(new_n267), .C2(new_n265), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n268), .B(new_n271), .C1(G77), .C2(new_n264), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n272), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT68), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n272), .A2(new_n283), .A3(new_n277), .A4(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G179), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(G20), .B1(new_n235), .B2(G50), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n232), .A2(new_n260), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n232), .A2(G33), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n288), .B1(new_n289), .B2(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n231), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n293), .A2(new_n295), .B1(new_n221), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n295), .B1(new_n273), .B2(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n221), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n282), .A2(new_n302), .A3(new_n284), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n287), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n282), .B2(new_n284), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n306), .A2(new_n307), .B1(new_n285), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n301), .B(KEYINPUT9), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n282), .A2(KEYINPUT72), .A3(G200), .A4(new_n284), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n309), .A2(new_n314), .A3(new_n310), .A4(new_n311), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n304), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n292), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n297), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n300), .B2(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(new_n295), .ZN(new_n320));
  XNOR2_X1  g0120(.A(G58), .B(G68), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G20), .A2(G33), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(G20), .B1(G159), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n261), .A2(new_n262), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n325), .A2(new_n326), .A3(G20), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n256), .A2(new_n257), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT7), .B1(new_n328), .B2(new_n232), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n330), .B2(G68), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n320), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n258), .A2(new_n263), .A3(new_n232), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n327), .B1(new_n326), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n323), .B1(new_n334), .B2(new_n210), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n319), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n325), .B1(G226), .B2(new_n265), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G223), .A2(G1698), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n279), .B1(new_n342), .B2(new_n271), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n275), .A2(new_n227), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT79), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G200), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n345), .A3(G190), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n338), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n338), .A2(KEYINPUT17), .A3(new_n347), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n338), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n346), .A2(new_n286), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n302), .B1(new_n343), .B2(new_n345), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(KEYINPUT18), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT80), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT18), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n356), .A2(new_n357), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n338), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n355), .A2(KEYINPUT80), .A3(KEYINPUT18), .A4(new_n358), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G238), .A2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n264), .B(new_n367), .C1(new_n227), .C2(G1698), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n271), .C1(G107), .C2(new_n264), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n280), .C1(new_n224), .C2(new_n275), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n286), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n292), .A2(new_n290), .B1(new_n232), .B2(new_n223), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT69), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n291), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n295), .B1(new_n223), .B2(new_n297), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n299), .A2(G77), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT70), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n370), .A2(new_n302), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n372), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n316), .A2(new_n354), .A3(new_n366), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n222), .A2(new_n265), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n227), .A2(G1698), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n264), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n270), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n279), .B1(new_n276), .B2(G238), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT13), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  INV_X1    g0192(.A(new_n387), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n258), .A2(new_n263), .B1(new_n227), .B2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n384), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n392), .B(new_n389), .C1(new_n395), .C2(new_n270), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT14), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n400), .A3(G169), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n391), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT73), .B(KEYINPUT13), .C1(new_n388), .C2(new_n390), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n386), .A2(new_n387), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n271), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT74), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n392), .A4(new_n389), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(G179), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT77), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n404), .A2(new_n405), .B1(new_n407), .B2(new_n411), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT77), .A3(G179), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n402), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n290), .B2(new_n221), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n210), .A2(G20), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n232), .A2(G33), .A3(G77), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n322), .A2(KEYINPUT75), .A3(G50), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n295), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT11), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT11), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n427), .A3(new_n295), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT12), .B1(new_n296), .B2(G68), .ZN(new_n431));
  AOI22_X1  g0231(.A1(G68), .A2(new_n299), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n429), .A2(KEYINPUT76), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT76), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n433), .A2(new_n434), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT78), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n418), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n416), .A2(G190), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n397), .A2(G200), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n435), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT71), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n377), .B2(new_n379), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n370), .A2(G200), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n448), .B1(new_n305), .B2(new_n370), .C1(new_n380), .C2(KEYINPUT71), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n442), .B(new_n445), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n383), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n273), .B(G45), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n455), .A2(new_n270), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G257), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n455), .A2(new_n278), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n256), .A2(new_n257), .A3(new_n255), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT67), .B1(new_n261), .B2(new_n262), .ZN(new_n462));
  OAI211_X1 g0262(.A(G250), .B(G1698), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G244), .B(new_n265), .C1(new_n256), .C2(new_n257), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n464), .A2(new_n465), .B1(G33), .B2(G283), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT81), .B1(new_n264), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT81), .ZN(new_n471));
  AOI211_X1 g0271(.A(new_n471), .B(new_n468), .C1(new_n258), .C2(new_n263), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n286), .B(new_n460), .C1(new_n473), .C2(new_n270), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT82), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n460), .B1(new_n473), .B2(new_n270), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n302), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n264), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n471), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n264), .A2(KEYINPUT81), .A3(new_n469), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(new_n466), .A3(new_n463), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n459), .B1(new_n481), .B2(new_n271), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n286), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n322), .A2(G77), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(KEYINPUT6), .A3(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n215), .A2(new_n486), .ZN(new_n488));
  NOR2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G20), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n485), .B(new_n492), .C1(new_n334), .C2(new_n486), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n295), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n273), .A2(G33), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n296), .A2(new_n495), .A3(new_n231), .A4(new_n294), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n215), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n296), .A2(G97), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n475), .A2(new_n477), .A3(new_n484), .A4(new_n501), .ZN(new_n502));
  AOI211_X1 g0302(.A(new_n497), .B(new_n499), .C1(new_n493), .C2(new_n295), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n482), .A2(G190), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n308), .C2(new_n482), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n213), .A2(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n264), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n513), .B(KEYINPUT22), .C1(new_n257), .C2(new_n256), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT86), .B1(new_n518), .B2(G20), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(new_n232), .A3(G33), .A4(G116), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n232), .B2(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n486), .A2(KEYINPUT23), .A3(G20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n517), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n512), .B1(new_n516), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT22), .B1(new_n264), .B2(new_n513), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n517), .A2(new_n522), .A3(new_n526), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n529), .A2(new_n511), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n510), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(KEYINPUT88), .A3(new_n295), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT88), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n511), .B1(new_n529), .B2(new_n530), .ZN(new_n535));
  INV_X1    g0335(.A(new_n513), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n258), .B2(new_n263), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n527), .B(new_n512), .C1(KEYINPUT22), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n509), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n534), .B1(new_n539), .B2(new_n320), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n214), .A2(new_n265), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n216), .A2(G1698), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n256), .C2(new_n257), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n271), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n455), .A2(G264), .A3(new_n270), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n458), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  INV_X1    g0350(.A(new_n549), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT25), .B1(new_n297), .B2(new_n486), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n486), .ZN(new_n555));
  INV_X1    g0355(.A(new_n496), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n554), .A2(new_n555), .B1(G107), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n541), .A2(new_n550), .A3(new_n552), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT88), .B1(new_n532), .B2(new_n295), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n539), .A2(new_n534), .A3(new_n320), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n551), .A2(G179), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT89), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n562), .B(new_n563), .C1(new_n302), .C2(new_n551), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n232), .B1(new_n387), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n489), .A2(new_n213), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n232), .B(G68), .C1(new_n256), .C2(new_n257), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n568), .B1(new_n291), .B2(new_n215), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n295), .ZN(new_n575));
  INV_X1    g0375(.A(new_n375), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n556), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n375), .A2(new_n297), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n211), .A2(new_n265), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n224), .A2(G1698), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n256), .C2(new_n257), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n518), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n271), .ZN(new_n584));
  INV_X1    g0384(.A(G45), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n214), .B1(new_n585), .B2(G1), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n273), .A2(new_n278), .A3(G45), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n270), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n286), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n270), .B1(new_n582), .B2(new_n518), .ZN(new_n590));
  INV_X1    g0390(.A(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n302), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n579), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n584), .A2(G190), .A3(new_n588), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n574), .A2(new_n295), .B1(new_n297), .B2(new_n375), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n556), .A2(G87), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT83), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT83), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n593), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n258), .A2(new_n263), .A3(G303), .ZN(new_n606));
  AND2_X1   g0406(.A1(G264), .A2(G1698), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n256), .B2(new_n257), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT84), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n325), .A2(KEYINPUT84), .A3(new_n607), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n325), .A2(G257), .A3(new_n265), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n606), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n271), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n456), .A2(G270), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n458), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G33), .A2(G283), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n232), .C1(G33), .C2(new_n215), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G20), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n295), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n294), .A2(new_n231), .B1(G20), .B2(new_n619), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(KEYINPUT20), .A3(new_n618), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n623), .A2(new_n625), .B1(G116), .B2(new_n556), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n297), .A2(new_n619), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n302), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n605), .B1(new_n616), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n614), .A2(G179), .A3(new_n458), .A4(new_n615), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n623), .A2(new_n625), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n556), .A2(G116), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n616), .A2(new_n628), .A3(new_n605), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n616), .A2(G200), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n638), .B(new_n634), .C1(new_n305), .C2(new_n616), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n603), .A2(new_n636), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n506), .A2(new_n558), .A3(new_n567), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n452), .A2(new_n641), .ZN(G372));
  NAND3_X1  g0442(.A1(new_n475), .A2(new_n477), .A3(new_n484), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n475), .A2(new_n477), .A3(new_n484), .A4(KEYINPUT90), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n599), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n501), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n593), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n506), .A2(new_n558), .A3(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n636), .A2(new_n637), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n565), .B1(new_n541), .B2(new_n557), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n564), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n502), .B1(new_n600), .B2(new_n602), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n651), .A2(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n451), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n359), .A2(new_n364), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n382), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n441), .B1(new_n662), .B2(new_n445), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n353), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n313), .A2(new_n315), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n304), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n666), .ZN(G369));
  INV_X1    g0467(.A(G13), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G20), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .A3(G1), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT27), .B1(new_n670), .B2(G1), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n634), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n652), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT91), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT91), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n677), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT92), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT92), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G330), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n561), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n558), .B1(new_n686), .B2(new_n676), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n567), .ZN(new_n688));
  INV_X1    g0488(.A(new_n567), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n676), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n675), .B1(new_n636), .B2(new_n637), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n567), .A2(new_n558), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n207), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n570), .A2(G116), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n699), .A2(new_n273), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n237), .B2(new_n699), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT28), .Z(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n656), .A2(new_n655), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n503), .B(new_n599), .C1(new_n645), .C2(new_n646), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n593), .B(new_n706), .C1(new_n707), .C2(new_n655), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT94), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n651), .A2(new_n654), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n649), .A2(KEYINPUT26), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT94), .A3(new_n593), .A4(new_n706), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n705), .B1(new_n714), .B2(new_n676), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n658), .A2(new_n705), .A3(new_n676), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n558), .A2(new_n502), .A3(new_n505), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n603), .A2(new_n636), .A3(new_n637), .A4(new_n639), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n564), .B2(new_n653), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n721), .A3(new_n676), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n547), .A2(new_n584), .A3(new_n548), .A4(new_n588), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n460), .B(new_n725), .C1(new_n473), .C2(new_n270), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n726), .B2(new_n630), .ZN(new_n727));
  INV_X1    g0527(.A(new_n630), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n482), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n584), .A2(new_n588), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n613), .A2(new_n271), .B1(G270), .B2(new_n456), .ZN(new_n731));
  AOI21_X1  g0531(.A(G179), .B1(new_n731), .B2(new_n458), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n476), .A2(new_n549), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n675), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n459), .B(new_n724), .C1(new_n481), .C2(new_n271), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT30), .B1(new_n736), .B2(new_n728), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n616), .A2(new_n286), .A3(new_n730), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n482), .A3(new_n551), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT93), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n727), .A2(new_n741), .A3(new_n733), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n729), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n675), .A2(KEYINPUT31), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n735), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n718), .B1(new_n722), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n715), .A2(new_n717), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n704), .B1(new_n747), .B2(G1), .ZN(G364));
  AOI21_X1  g0548(.A(new_n273), .B1(new_n669), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n699), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(G355), .A2(new_n207), .A3(new_n264), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n698), .A2(new_n325), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n236), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n250), .A2(new_n585), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n752), .B1(G116), .B2(new_n207), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n231), .B1(G20), .B2(new_n302), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n232), .A2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n264), .B1(G329), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n232), .A2(new_n305), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n286), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n769), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n286), .A2(new_n308), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G326), .ZN(new_n778));
  INV_X1    g0578(.A(G294), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n766), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n765), .A2(new_n772), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n778), .B1(new_n779), .B2(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT98), .Z(new_n786));
  INV_X1    g0586(.A(G317), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT33), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(new_n765), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(KEYINPUT33), .B2(new_n787), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n774), .B(new_n786), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n765), .A2(new_n286), .A3(G200), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n771), .A2(new_n286), .A3(G200), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n791), .B1(new_n792), .B2(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n776), .A2(new_n221), .B1(new_n784), .B2(new_n223), .ZN(new_n800));
  INV_X1    g0600(.A(new_n773), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G58), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n781), .A2(G97), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n796), .A2(new_n486), .B1(new_n210), .B2(new_n789), .ZN(new_n806));
  INV_X1    g0606(.A(new_n798), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G87), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n767), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n264), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n799), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n762), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n751), .B(new_n764), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n683), .A2(new_n684), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n761), .ZN(new_n817));
  INV_X1    g0617(.A(new_n685), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n751), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n718), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n658), .A2(new_n676), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n382), .A2(new_n675), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n380), .A2(new_n675), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n449), .B2(new_n447), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n824), .B1(new_n826), .B2(new_n382), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n676), .B(new_n827), .C1(new_n650), .C2(new_n657), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(new_n746), .ZN(new_n832));
  INV_X1    g0632(.A(new_n751), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n264), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n835), .B1(new_n797), .B2(new_n776), .C1(new_n783), .C2(new_n767), .ZN(new_n836));
  INV_X1    g0636(.A(new_n796), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G87), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n801), .A2(G294), .ZN(new_n839));
  INV_X1    g0639(.A(new_n784), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G116), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n804), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n836), .B(new_n842), .C1(G107), .C2(new_n807), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n792), .B2(new_n789), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n837), .A2(G68), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n221), .B2(new_n798), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n328), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n226), .B2(new_n782), .C1(new_n850), .C2(new_n767), .ZN(new_n851));
  INV_X1    g0651(.A(new_n789), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G143), .A2(new_n801), .B1(new_n852), .B2(G150), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n777), .A2(G137), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n809), .C2(new_n784), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT34), .Z(new_n856));
  OAI21_X1  g0656(.A(new_n845), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT102), .Z(new_n858));
  AOI21_X1  g0658(.A(new_n833), .B1(new_n858), .B2(new_n762), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n762), .A2(new_n757), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT99), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n223), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n859), .B(new_n862), .C1(new_n758), .C2(new_n827), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n834), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NAND2_X1  g0665(.A1(new_n366), .A2(new_n354), .ZN(new_n866));
  INV_X1    g0666(.A(new_n673), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n332), .B1(KEYINPUT16), .B2(new_n331), .ZN(new_n868));
  INV_X1    g0668(.A(new_n319), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n349), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n338), .B1(new_n363), .B2(new_n673), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT37), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n363), .A2(new_n673), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n870), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(new_n349), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n355), .B(new_n867), .C1(new_n660), .C2(new_n353), .ZN(new_n882));
  INV_X1    g0682(.A(new_n873), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n875), .A3(new_n349), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n872), .B2(new_n873), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(KEYINPUT37), .C1(new_n872), .C2(new_n873), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n881), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n871), .A2(new_n880), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n890), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n442), .A2(new_n675), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n824), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n830), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n436), .A2(new_n439), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n399), .A2(new_n401), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n413), .A2(new_n414), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT77), .B1(new_n416), .B2(G179), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n445), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n902), .B(new_n675), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n675), .B1(new_n436), .B2(new_n439), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n445), .B(new_n909), .C1(new_n418), .C2(new_n440), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n871), .B2(new_n880), .ZN(new_n912));
  INV_X1    g0712(.A(new_n870), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n366), .B2(new_n354), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n890), .B(new_n879), .C1(new_n914), .C2(new_n867), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n901), .B(new_n911), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n660), .A2(new_n673), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n899), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT105), .Z(new_n919));
  OAI21_X1  g0719(.A(new_n451), .B1(new_n715), .B2(new_n717), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n666), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n915), .A2(new_n912), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n828), .B1(new_n910), .B2(new_n908), .ZN(new_n925));
  INV_X1    g0725(.A(new_n735), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n734), .A2(new_n744), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n926), .B(new_n927), .C1(new_n641), .C2(new_n675), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n923), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n925), .A4(new_n928), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(G330), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(G330), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n452), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(new_n928), .A3(new_n931), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n934), .B1(new_n452), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n922), .B(new_n936), .Z(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n273), .B2(new_n669), .ZN(new_n938));
  OAI21_X1  g0738(.A(G77), .B1(new_n226), .B2(new_n210), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n236), .A2(new_n939), .B1(G50), .B2(new_n210), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n668), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n619), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n233), .C1(KEYINPUT35), .C2(new_n491), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n941), .A3(new_n945), .ZN(G367));
  AOI22_X1  g0746(.A1(G311), .A2(new_n777), .B1(new_n801), .B2(G303), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n947), .B(new_n328), .C1(new_n787), .C2(new_n767), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G283), .B2(new_n840), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n798), .A2(new_n619), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT46), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G107), .B2(new_n781), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n837), .A2(G97), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n852), .A2(G294), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n949), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n840), .A2(G50), .B1(new_n781), .B2(G68), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n809), .B2(new_n789), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G137), .B2(new_n768), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n837), .A2(G77), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n777), .A2(G143), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n264), .B1(new_n289), .B2(new_n773), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G58), .B2(new_n807), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT107), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n833), .B1(new_n966), .B2(new_n762), .ZN(new_n967));
  INV_X1    g0767(.A(new_n753), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n763), .B1(new_n207), .B2(new_n375), .C1(new_n241), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n596), .A2(new_n597), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n675), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n648), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n593), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n967), .B(new_n969), .C1(new_n760), .C2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n506), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n695), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n979));
  INV_X1    g0779(.A(new_n502), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n647), .A2(new_n501), .A3(new_n675), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n506), .B1(new_n503), .B2(new_n676), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n980), .B1(new_n983), .B2(new_n689), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n979), .B1(new_n984), .B2(new_n675), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT106), .Z(new_n986));
  OR2_X1    g0786(.A1(new_n978), .A2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT43), .ZN(new_n993));
  INV_X1    g0793(.A(new_n974), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n986), .A2(new_n993), .A3(new_n994), .A4(new_n987), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n692), .A2(new_n983), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n992), .A2(new_n692), .A3(new_n983), .A4(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n696), .A2(new_n983), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT45), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n696), .A2(new_n983), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n692), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n694), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n691), .A2(new_n1007), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n685), .A2(new_n1008), .A3(new_n695), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n685), .B1(new_n1008), .B2(new_n695), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n747), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n699), .B(KEYINPUT41), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n750), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n975), .B1(new_n1000), .B2(new_n1014), .ZN(G387));
  NAND3_X1  g0815(.A1(new_n701), .A2(new_n207), .A3(new_n264), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n246), .A2(G45), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n968), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n292), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  AOI21_X1  g0819(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT50), .B1(new_n292), .B2(G50), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1019), .A2(new_n700), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1018), .A2(new_n1022), .B1(new_n486), .B2(new_n698), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n763), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n751), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT108), .B(G322), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n777), .A2(new_n1026), .B1(new_n801), .B2(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n797), .B2(new_n784), .C1(new_n783), .C2(new_n789), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n792), .B2(new_n782), .C1(new_n779), .C2(new_n798), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT49), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n325), .B1(new_n768), .B2(G326), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n619), .C2(new_n796), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n325), .B1(new_n784), .B2(new_n210), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n576), .A2(new_n781), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n807), .A2(G77), .B1(new_n801), .B2(G50), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n953), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1034), .B(new_n1037), .C1(G150), .C2(new_n768), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n809), .B2(new_n776), .C1(new_n292), .C2(new_n789), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n814), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1025), .B(new_n1040), .C1(new_n691), .C2(new_n761), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1011), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n750), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n747), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n699), .B1(new_n1042), .B2(new_n747), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(G393));
  XNOR2_X1  g0847(.A(new_n1005), .B(new_n693), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n699), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1006), .B2(new_n1044), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1048), .A2(new_n750), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n835), .B1(new_n779), .B2(new_n784), .C1(new_n797), .C2(new_n789), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n776), .A2(new_n787), .B1(new_n773), .B2(new_n783), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT52), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n486), .B2(new_n796), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1054), .B(new_n1057), .C1(G116), .C2(new_n781), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n768), .A2(new_n1026), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n792), .C2(new_n798), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT109), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n776), .A2(new_n289), .B1(new_n773), .B2(new_n809), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT51), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1062), .A2(new_n1063), .B1(G77), .B2(new_n781), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n840), .A2(new_n317), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n838), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n798), .A2(new_n210), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n768), .A2(G143), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n325), .B1(new_n789), .B2(new_n221), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n762), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n763), .B1(new_n215), .B2(new_n207), .C1(new_n253), .C2(new_n968), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n981), .A2(new_n982), .A3(new_n761), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1072), .A2(new_n751), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1052), .A2(new_n1053), .A3(new_n1075), .ZN(G390));
  NAND2_X1  g0876(.A1(new_n901), .A2(new_n911), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n898), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n894), .A2(new_n897), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n746), .A2(new_n827), .A3(new_n911), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n911), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n826), .A2(new_n382), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n714), .A2(new_n676), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n1085), .B2(new_n900), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n892), .A2(new_n1078), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1081), .B(new_n1082), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n900), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n911), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1087), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1090), .A2(new_n1091), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n911), .A2(new_n928), .A3(G330), .A4(new_n827), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n928), .A2(G330), .A3(new_n827), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1083), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1096), .A2(new_n1082), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1097), .A2(new_n900), .A3(new_n1085), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n911), .B1(new_n746), .B2(new_n827), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT111), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(KEYINPUT111), .B(new_n911), .C1(new_n746), .C2(new_n827), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n901), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT112), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT112), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n901), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT110), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n452), .B2(new_n933), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n933), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n451), .A2(KEYINPUT110), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n920), .A3(new_n666), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1094), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1081), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n925), .A3(new_n1110), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1088), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1118), .A3(new_n699), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1094), .A2(new_n749), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1080), .A2(new_n757), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n789), .A2(new_n486), .B1(new_n784), .B2(new_n215), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT113), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n792), .C2(new_n776), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT114), .Z(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n264), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n801), .A2(G116), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n807), .A2(G87), .B1(G77), .B2(new_n781), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n846), .B1(new_n779), .B2(new_n767), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT115), .Z(new_n1132));
  NAND4_X1  g0932(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n837), .A2(G50), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n798), .A2(new_n289), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n852), .A2(G137), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n777), .B1(new_n801), .B2(G132), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  AOI211_X1 g0940(.A(new_n835), .B(new_n1139), .C1(new_n840), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n768), .A2(G125), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n809), .C2(new_n782), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n814), .B1(new_n1133), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n833), .B(new_n1144), .C1(new_n292), .C2(new_n861), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1121), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1120), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1119), .A2(new_n1147), .ZN(G378));
  XOR2_X1   g0948(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n316), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n301), .A2(new_n867), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n316), .A2(new_n1150), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n932), .A2(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1160), .A2(new_n930), .A3(G330), .A4(new_n931), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1159), .A2(new_n918), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n918), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n750), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n782), .A2(new_n210), .B1(new_n776), .B2(new_n619), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT116), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n837), .A2(G58), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n798), .A2(new_n223), .B1(new_n789), .B2(new_n215), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G41), .B(new_n1169), .C1(new_n576), .C2(new_n840), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n328), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n486), .B2(new_n773), .C1(new_n792), .C2(new_n767), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(G124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n260), .B1(new_n767), .B2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G128), .A2(new_n801), .B1(new_n840), .B2(G137), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n807), .A2(new_n1140), .B1(G150), .B2(new_n781), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n852), .A2(G132), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n777), .A2(G125), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1182));
  AOI211_X1 g0982(.A(G41), .B(new_n1176), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n809), .B2(new_n796), .C1(new_n1182), .C2(new_n1181), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n221), .B1(new_n256), .B2(G41), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n762), .B1(new_n1174), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT119), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n833), .B1(new_n221), .B2(new_n860), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(new_n1158), .C2(new_n758), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1165), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1113), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1094), .B2(new_n1107), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(KEYINPUT57), .A3(new_n1164), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n699), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1164), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1191), .B1(new_n1195), .B2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n852), .A2(new_n1140), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1168), .B(new_n1198), .C1(new_n221), .C2(new_n782), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n328), .B(new_n1199), .C1(G150), .C2(new_n840), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G137), .A2(new_n801), .B1(new_n768), .B2(G128), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n850), .B2(new_n776), .C1(new_n809), .C2(new_n798), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n959), .B1(new_n779), .B2(new_n776), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n789), .A2(new_n619), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1035), .B1(new_n486), .B2(new_n784), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n835), .B1(new_n215), .B2(new_n798), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n792), .B2(new_n773), .C1(new_n797), .C2(new_n767), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n814), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n833), .B(new_n1210), .C1(new_n210), .C2(new_n861), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n758), .B2(new_n911), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1107), .B2(new_n749), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1013), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n1216), .B2(new_n1115), .ZN(G381));
  NOR2_X1   g1017(.A1(G375), .A2(G378), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(G384), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT120), .Z(new_n1222));
  AND3_X1   g1022(.A1(new_n1052), .A2(new_n1053), .A3(new_n1075), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n975), .C1(new_n1014), .C2(new_n1000), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G381), .A2(new_n1219), .A3(new_n1222), .A4(new_n1224), .ZN(G407));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G343), .C2(new_n1219), .ZN(G409));
  OAI21_X1  g1026(.A(KEYINPUT60), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1215), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1113), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n699), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1228), .A2(KEYINPUT121), .A3(new_n699), .A4(new_n1229), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1214), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n864), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(G384), .A3(new_n1214), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1238), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G384), .B1(new_n1234), .B2(new_n1214), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n864), .B(new_n1213), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1191), .B(G378), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1193), .A2(new_n1013), .A3(new_n1164), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1165), .A2(new_n1190), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1147), .B(new_n1119), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n674), .A2(G213), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1239), .A2(new_n1243), .A3(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1236), .A3(new_n1237), .A4(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT63), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(G390), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1224), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT122), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1220), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1262), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1260), .B1(new_n1220), .B2(new_n1261), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1224), .B(new_n1258), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1257), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(KEYINPUT123), .B(KEYINPUT61), .C1(new_n1263), .C2(new_n1266), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1254), .A2(new_n1256), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT124), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1263), .A2(new_n1273), .A3(new_n1266), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1252), .A2(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1268), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1272), .A2(new_n1280), .ZN(G405));
  NAND3_X1  g1081(.A1(G375), .A2(new_n1147), .A3(new_n1119), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT125), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1241), .A2(new_n1242), .A3(KEYINPUT125), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1244), .B(new_n1282), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1284), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1244), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1276), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT126), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1267), .A2(KEYINPUT124), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1263), .A2(new_n1273), .A3(new_n1266), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1291), .A3(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1296), .A3(new_n1289), .A4(new_n1286), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1292), .A2(new_n1297), .ZN(G402));
endmodule


