//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT91), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G122), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT83), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(new_n192), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT67), .A2(G116), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n193), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT5), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n197), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n195), .A2(G119), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n193), .A2(KEYINPUT66), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n202), .B(G116), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G113), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT81), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(G116), .B1(new_n204), .B2(new_n205), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n200), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT67), .A2(G116), .ZN(new_n213));
  OAI21_X1  g027(.A(G119), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(G107), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n216), .B(new_n219), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n209), .A2(KEYINPUT5), .A3(new_n214), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G113), .A4(new_n206), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n208), .A2(new_n215), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n210), .B1(new_n197), .B2(new_n201), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n215), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n237), .A3(G101), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n231), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n231), .B2(new_n239), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT6), .B(new_n191), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n231), .A2(new_n239), .A3(new_n190), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT84), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n231), .A2(new_n239), .A3(new_n248), .A4(new_n190), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n191), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n231), .A2(new_n239), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n253), .B2(new_n241), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n244), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  OAI211_X1 g074(.A(G128), .B(new_n257), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n262), .B(new_n263), .C1(KEYINPUT1), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT75), .A2(G125), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT75), .A2(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n269), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n262), .A2(new_n263), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT64), .ZN(new_n277));
  XNOR2_X1  g091(.A(G143), .B(G146), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n273), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n277), .A2(new_n262), .A3(new_n263), .A4(new_n273), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n270), .B1(new_n271), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G224), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n284), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n255), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT87), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n255), .A2(new_n287), .A3(KEYINPUT87), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n262), .A2(new_n263), .A3(new_n273), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT64), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n278), .A2(new_n277), .A3(new_n273), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n294), .A2(new_n295), .B1(new_n272), .B2(new_n275), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n270), .A2(KEYINPUT88), .B1(new_n269), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n270), .A2(KEYINPUT88), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n299));
  OAI22_X1  g113(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n286), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT89), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n300), .A2(KEYINPUT89), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n286), .B2(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n282), .B(new_n304), .C1(new_n303), .C2(new_n286), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n190), .B(KEYINPUT8), .Z(new_n306));
  OAI21_X1  g120(.A(new_n215), .B1(new_n203), .B2(new_n207), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(new_n227), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n208), .A2(new_n215), .A3(new_n230), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(new_n227), .ZN(new_n310));
  AND4_X1   g124(.A1(new_n301), .A2(new_n302), .A3(new_n305), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n247), .A2(new_n249), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n189), .B1(new_n292), .B2(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n255), .A2(new_n287), .A3(KEYINPUT87), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT87), .B1(new_n255), .B2(new_n287), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n189), .B(new_n313), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G214), .B1(G237), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(G234), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n267), .A2(G140), .A3(new_n268), .ZN(new_n328));
  OR2_X1    g142(.A1(G125), .A2(G140), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(KEYINPUT16), .A2(G140), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n269), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G146), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n259), .B1(new_n330), .B2(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n264), .B1(new_n194), .B2(new_n196), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n193), .A2(G128), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(KEYINPUT23), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n204), .A2(new_n205), .A3(G128), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(KEYINPUT23), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G110), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT72), .B1(new_n337), .B2(new_n338), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT72), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT66), .B(G119), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(new_n264), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n346), .B2(new_n350), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT24), .B(G110), .Z(new_n355));
  AOI21_X1  g169(.A(new_n345), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n350), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n355), .A3(new_n351), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n344), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n355), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n352), .B2(new_n353), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n341), .A2(G110), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n334), .A2(KEYINPUT76), .ZN(new_n366));
  NOR4_X1   g180(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT76), .A4(new_n259), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n259), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT22), .B(G137), .ZN(new_n373));
  INV_X1    g187(.A(G221), .ZN(new_n374));
  INV_X1    g188(.A(G234), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(G953), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n373), .B(new_n376), .Z(new_n377));
  NAND3_X1  g191(.A1(new_n361), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n354), .A2(new_n345), .A3(new_n355), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n343), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n333), .B2(G146), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n371), .B1(new_n384), .B2(new_n367), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n364), .B2(new_n363), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n387), .A3(new_n324), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n378), .A2(new_n387), .A3(KEYINPUT25), .A4(new_n324), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n326), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n325), .A2(G902), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n378), .A2(new_n387), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n398));
  INV_X1    g212(.A(G134), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(G137), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(G137), .ZN(new_n401));
  INV_X1    g215(.A(G137), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT65), .A3(G134), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G131), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT11), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n399), .B2(G137), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(KEYINPUT11), .A3(G134), .ZN(new_n408));
  INV_X1    g222(.A(G131), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n401), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n405), .A2(new_n410), .A3(new_n265), .A4(new_n261), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n408), .A3(new_n401), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G131), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(new_n414), .B2(new_n281), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n233), .ZN(new_n416));
  INV_X1    g230(.A(new_n233), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n410), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n296), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n419), .A3(new_n411), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(KEYINPUT69), .A3(new_n420), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n415), .A2(KEYINPUT69), .A3(new_n233), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT28), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n421), .A2(new_n422), .A3(new_n426), .A4(KEYINPUT28), .ZN(new_n429));
  INV_X1    g243(.A(G237), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n285), .A3(G210), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(G101), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(KEYINPUT29), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT71), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n415), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n233), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n420), .ZN(new_n442));
  INV_X1    g256(.A(new_n434), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(KEYINPUT68), .A3(new_n443), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT28), .A4(new_n411), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n425), .A2(new_n448), .A3(new_n416), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT29), .B1(new_n449), .B2(new_n434), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n428), .A2(new_n452), .A3(new_n429), .A4(new_n435), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n437), .A2(new_n451), .A3(new_n324), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G472), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n441), .A2(new_n434), .A3(new_n420), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT31), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT31), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n441), .A2(new_n458), .A3(new_n434), .A4(new_n420), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n457), .B(new_n459), .C1(new_n434), .C2(new_n449), .ZN(new_n460));
  NOR2_X1   g274(.A1(G472), .A2(G902), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n460), .A2(KEYINPUT32), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT32), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n397), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n264), .A2(G143), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n399), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n256), .A2(G128), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n469), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G122), .B1(new_n212), .B2(new_n213), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n192), .B2(G122), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n476), .A2(G107), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(G107), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n192), .A2(G122), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n475), .B2(KEYINPUT14), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n481), .A2(KEYINPUT94), .B1(KEYINPUT14), .B2(new_n475), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n481), .A2(KEYINPUT94), .ZN(new_n483));
  OAI21_X1  g297(.A(G107), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n473), .B(G134), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n479), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT9), .B(G234), .Z(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(G217), .A3(new_n285), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n487), .B(new_n489), .Z(new_n490));
  AOI211_X1 g304(.A(KEYINPUT15), .B(new_n468), .C1(new_n490), .C2(new_n324), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n324), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n430), .A2(new_n285), .A3(G214), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(G143), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n409), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT18), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n497), .B1(new_n500), .B2(new_n409), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n328), .A2(G146), .A3(new_n329), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n371), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(KEYINPUT17), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n496), .B(new_n256), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G131), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n497), .A2(new_n409), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n505), .B1(new_n509), .B2(KEYINPUT17), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n504), .B1(new_n510), .B2(new_n336), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n220), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n511), .A2(new_n514), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n324), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G475), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n384), .A2(new_n367), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n328), .A2(KEYINPUT19), .A3(new_n329), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT19), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n370), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT92), .B1(new_n523), .B2(G146), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n520), .A2(new_n525), .A3(new_n259), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n509), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n504), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n513), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT93), .B(new_n504), .C1(new_n519), .C2(new_n527), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G475), .A2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT20), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n532), .A2(KEYINPUT20), .A3(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n518), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n495), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n374), .B1(new_n488), .B2(new_n324), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n236), .A2(new_n296), .A3(new_n238), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n261), .A2(new_n265), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n227), .A2(new_n542), .A3(KEYINPUT10), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n223), .A2(new_n261), .A3(new_n265), .A4(new_n225), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT10), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n541), .A2(new_n543), .A3(new_n414), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n226), .A2(new_n266), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n544), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n549), .A2(KEYINPUT12), .A3(new_n418), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT12), .B1(new_n549), .B2(new_n418), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n285), .A2(G227), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT78), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G140), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n547), .A2(new_n556), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n541), .A2(new_n546), .A3(new_n543), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n418), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n552), .A2(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT79), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n324), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G469), .ZN(new_n565));
  INV_X1    g379(.A(G469), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n547), .B(new_n556), .C1(new_n550), .C2(new_n551), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n556), .B1(new_n560), .B2(new_n547), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n566), .B(new_n324), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT80), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n560), .A2(new_n547), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n557), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n567), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(KEYINPUT80), .A3(new_n566), .A4(new_n324), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n540), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n285), .A2(G952), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n375), .B2(new_n430), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n324), .B(new_n285), .C1(G234), .C2(G237), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT21), .B(G898), .Z(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n539), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n322), .A2(new_n467), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  AOI21_X1  g401(.A(new_n321), .B1(new_n314), .B2(KEYINPUT95), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n188), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n317), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n487), .B(new_n489), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n594), .A2(KEYINPUT33), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(KEYINPUT33), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(G478), .A3(new_n324), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n492), .A2(new_n468), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n532), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT20), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n533), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n603), .A2(new_n535), .B1(G475), .B2(new_n517), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n584), .ZN(new_n606));
  INV_X1    g420(.A(G472), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n460), .B2(new_n324), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n460), .B2(new_n461), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n397), .A2(new_n578), .A3(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n593), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND3_X1  g427(.A1(new_n495), .A2(new_n584), .A3(new_n604), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n593), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT96), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NAND2_X1  g432(.A1(new_n390), .A2(new_n391), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n325), .ZN(new_n620));
  OAI22_X1  g434(.A1(new_n382), .A2(new_n386), .B1(KEYINPUT36), .B2(new_n379), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n379), .A2(KEYINPUT36), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n361), .A2(new_n372), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n394), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n322), .A2(new_n585), .A3(new_n609), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  AND3_X1   g443(.A1(new_n465), .A2(new_n578), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n495), .A2(new_n604), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n581), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n580), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n630), .A2(new_n588), .A3(new_n592), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  INV_X1    g452(.A(new_n464), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n421), .A2(new_n422), .A3(new_n443), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n456), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n607), .B1(new_n641), .B2(new_n324), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n643), .A2(new_n321), .A3(new_n626), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n495), .A3(new_n538), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n590), .A2(new_n317), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n634), .B(KEYINPUT39), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n578), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT40), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n645), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT98), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n256), .ZN(G45));
  NAND3_X1  g469(.A1(new_n538), .A2(new_n599), .A3(new_n634), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n630), .A2(new_n588), .A3(new_n592), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  AOI21_X1  g473(.A(new_n566), .B1(new_n575), .B2(new_n324), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT99), .ZN(new_n661));
  INV_X1    g475(.A(new_n540), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n661), .A2(new_n662), .A3(new_n577), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n593), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n467), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n606), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT41), .B(G113), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G15));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n614), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n192), .ZN(G18));
  AND4_X1   g485(.A1(new_n465), .A2(new_n539), .A3(new_n584), .A4(new_n626), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT100), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n193), .ZN(G21));
  INV_X1    g489(.A(new_n665), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n495), .A2(new_n538), .A3(KEYINPUT101), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n491), .A2(new_n494), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n604), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n428), .A2(new_n429), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n457), .B(new_n459), .C1(new_n682), .C2(new_n434), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n608), .B1(new_n683), .B2(new_n461), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n397), .A3(new_n584), .A4(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n676), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(G122), .Z(G24));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n461), .ZN(new_n688));
  INV_X1    g502(.A(new_n608), .ZN(new_n689));
  INV_X1    g503(.A(new_n625), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n688), .B(new_n689), .C1(new_n392), .C2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n656), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n588), .A2(new_n692), .A3(new_n592), .A4(new_n663), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  NOR2_X1   g508(.A1(new_n646), .A2(new_n321), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n561), .B2(G902), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n540), .B1(new_n577), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n695), .A2(new_n467), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n656), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G131), .ZN(G33));
  NAND4_X1  g519(.A1(new_n695), .A2(new_n467), .A3(new_n636), .A4(new_n697), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  NOR2_X1   g521(.A1(new_n600), .A2(new_n538), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT43), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT103), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT103), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n392), .A2(new_n690), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n609), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n562), .A2(new_n718), .A3(new_n563), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n566), .B1(new_n561), .B2(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(G469), .A2(G902), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT46), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n724), .A2(KEYINPUT46), .B1(new_n572), .B2(new_n576), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n540), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n650), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n716), .A2(new_n695), .A3(new_n717), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G137), .ZN(G39));
  NOR2_X1   g545(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n732));
  AND2_X1   g546(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n727), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n727), .B2(new_n732), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n656), .A2(new_n397), .A3(new_n465), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n695), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G140), .ZN(G42));
  INV_X1    g553(.A(new_n643), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n661), .A2(new_n577), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n740), .B1(KEYINPUT49), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n742), .A2(KEYINPUT49), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n397), .A2(new_n708), .A3(new_n320), .A4(new_n662), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n648), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n637), .A2(new_n658), .A3(new_n693), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n620), .A2(new_n697), .A3(new_n625), .A4(new_n634), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n392), .A2(new_n690), .A3(new_n635), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n697), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n740), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n588), .A2(new_n681), .A3(new_n592), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n748), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n748), .B2(new_n756), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n589), .A2(KEYINPUT95), .A3(new_n188), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n320), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n319), .B2(new_n591), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n764), .B(new_n630), .C1(new_n636), .C2(new_n657), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n712), .A2(new_n751), .A3(new_n634), .A4(new_n697), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n643), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n764), .A2(new_n768), .A3(new_n681), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(KEYINPUT107), .A3(new_n693), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(new_n761), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n759), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g587(.A(KEYINPUT108), .B(KEYINPUT52), .C1(new_n761), .C2(new_n770), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT109), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n637), .A2(new_n658), .A3(new_n693), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT107), .B1(new_n776), .B2(new_n769), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n748), .A2(new_n756), .A3(new_n760), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n757), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n771), .A2(new_n772), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n759), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n674), .ZN(new_n785));
  OAI22_X1  g599(.A1(new_n666), .A2(new_n606), .B1(new_n676), .B2(new_n685), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n670), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n610), .B1(new_n606), .B2(new_n614), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n322), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n627), .A2(new_n789), .A3(new_n586), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n695), .A2(new_n539), .A3(new_n634), .A4(new_n630), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n695), .A2(new_n692), .A3(new_n697), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n706), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n785), .A2(new_n704), .A3(new_n787), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT53), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n761), .A2(new_n770), .A3(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n779), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n674), .A2(new_n670), .A3(new_n786), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT112), .B1(new_n790), .B2(new_n793), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(new_n704), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n775), .B2(new_n783), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n800), .B1(new_n795), .B2(new_n798), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n804), .B1(new_n803), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n580), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n397), .A2(new_n709), .A3(new_n818), .A4(new_n684), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n321), .A3(new_n648), .A4(new_n663), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT50), .Z(new_n821));
  NOR4_X1   g635(.A1(new_n664), .A2(new_n646), .A3(new_n321), .A4(new_n580), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n397), .A3(new_n643), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT114), .Z(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n604), .A3(new_n600), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n822), .A2(new_n709), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n626), .A3(new_n684), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT51), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n735), .B1(new_n662), .B2(new_n742), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n695), .A3(new_n819), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n829), .B(new_n833), .C1(new_n830), .C2(KEYINPUT51), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n826), .A2(new_n467), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n819), .A2(new_n665), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n579), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n605), .B2(new_n824), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n835), .A2(new_n836), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n805), .A2(new_n817), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(G952), .A2(G953), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT115), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n747), .B1(new_n844), .B2(new_n846), .ZN(G75));
  INV_X1    g661(.A(new_n811), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n758), .B1(new_n779), .B2(KEYINPUT108), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n781), .B1(new_n849), .B2(new_n782), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n773), .A2(KEYINPUT109), .A3(new_n774), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n799), .A2(new_n801), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(G902), .A3(new_n188), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n255), .B(new_n287), .Z(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT55), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(KEYINPUT117), .A3(new_n859), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n285), .A2(G952), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n855), .B2(KEYINPUT116), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n857), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n869), .ZN(G51));
  XNOR2_X1  g684(.A(new_n814), .B(KEYINPUT54), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n722), .B(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n575), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n814), .A2(new_n324), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n719), .A3(new_n720), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n864), .B1(new_n873), .B2(new_n875), .ZN(G54));
  NAND3_X1  g690(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT118), .B1(new_n877), .B2(new_n532), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n864), .B1(new_n877), .B2(new_n532), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n532), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(G60));
  AND2_X1   g696(.A1(new_n595), .A2(new_n596), .ZN(new_n883));
  NAND2_X1  g697(.A1(G478), .A2(G902), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT59), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n865), .B1(new_n871), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n805), .B2(new_n817), .ZN(new_n888));
  INV_X1    g702(.A(new_n883), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G63));
  XNOR2_X1  g704(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n323), .A2(new_n324), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n812), .B2(new_n813), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n864), .B1(new_n894), .B2(new_n395), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n624), .B(new_n893), .C1(new_n812), .C2(new_n813), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(KEYINPUT61), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n854), .A2(new_n898), .A3(new_n624), .A4(new_n893), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n895), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(G66));
  AOI21_X1  g720(.A(new_n285), .B1(new_n583), .B2(G224), .ZN(new_n907));
  INV_X1    g721(.A(new_n790), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n806), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT122), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(new_n910), .B2(new_n285), .ZN(new_n911));
  INV_X1    g725(.A(new_n255), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(G898), .B2(new_n285), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n911), .B(new_n913), .Z(G69));
  INV_X1    g728(.A(G227), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n915), .B2(new_n632), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n439), .A2(new_n440), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT123), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n523), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT125), .B(G900), .Z(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT126), .Z(new_n922));
  NOR2_X1   g736(.A1(new_n654), .A2(new_n748), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(KEYINPUT124), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n730), .A2(new_n738), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n923), .A2(KEYINPUT124), .A3(new_n924), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n466), .A2(new_n651), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n631), .B1(new_n604), .B2(new_n600), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n695), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n927), .A2(new_n929), .A3(new_n930), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n919), .B1(new_n934), .B2(new_n285), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n729), .A2(new_n467), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n704), .B(new_n706), .C1(new_n755), .C2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n928), .A2(new_n937), .A3(new_n748), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n919), .A2(new_n285), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n916), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n922), .B1(new_n935), .B2(new_n940), .ZN(G72));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT63), .Z(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n934), .B2(new_n910), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n434), .A3(new_n442), .ZN(new_n945));
  INV_X1    g759(.A(new_n938), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n946), .B2(new_n910), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n442), .A2(new_n434), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT127), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n864), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n796), .A2(new_n802), .ZN(new_n952));
  INV_X1    g766(.A(new_n943), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n446), .A2(new_n447), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n456), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n952), .B2(new_n955), .ZN(G57));
endmodule


