//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n205), .A2(new_n207), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n213), .A2(new_n214), .A3(new_n208), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n213), .A2(new_n208), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n218));
  AND2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(new_n206), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT24), .A3(new_n212), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n218), .A2(new_n221), .A3(KEYINPUT25), .A4(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT26), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n231), .B(new_n212), .C1(new_n233), .C2(new_n219), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G183gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n237), .A3(new_n223), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n234), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT66), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n234), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .A4(new_n223), .ZN(new_n250));
  AND4_X1   g049(.A1(KEYINPUT66), .A2(new_n246), .A3(new_n244), .A4(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n228), .B(new_n230), .C1(new_n245), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT1), .B1(new_n253), .B2(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(G134gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G127gat), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G113gat), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n254), .B(new_n256), .C1(KEYINPUT69), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G120gat), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n261), .A2(new_n258), .A3(KEYINPUT69), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT1), .B1(new_n261), .B2(new_n258), .ZN(new_n264));
  OR2_X1    g063(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(G127gat), .A3(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n255), .A2(G127gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(KEYINPUT68), .A3(new_n269), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n244), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n246), .A2(new_n244), .A3(new_n250), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n281), .A2(new_n282), .A3(new_n253), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n271), .B1(new_n283), .B2(new_n268), .ZN(new_n284));
  INV_X1    g083(.A(new_n264), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n273), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n263), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n280), .A2(new_n288), .A3(new_n228), .A4(new_n230), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n275), .A2(new_n289), .B1(G227gat), .B2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT34), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT34), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT72), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n289), .ZN(new_n296));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n290), .A2(new_n300), .A3(new_n294), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n293), .A2(new_n295), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n275), .A2(G227gat), .A3(G233gat), .A4(new_n289), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n304));
  XNOR2_X1  g103(.A(G15gat), .B(G43gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT70), .ZN(new_n306));
  XNOR2_X1  g105(.A(G71gat), .B(G99gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n303), .B(KEYINPUT32), .C1(new_n304), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT33), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n303), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314));
  AOI211_X1 g113(.A(new_n314), .B(new_n308), .C1(new_n303), .C2(new_n311), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n302), .B(new_n309), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n309), .B1(new_n313), .B2(new_n315), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n295), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n301), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324));
  INV_X1    g123(.A(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G141gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n326), .A2(new_n328), .B1(KEYINPUT2), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n329), .ZN(new_n335));
  AND2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT78), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(new_n337), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(KEYINPUT77), .ZN(new_n342));
  XNOR2_X1  g141(.A(G141gat), .B(G148gat), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n324), .B1(new_n274), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n346), .A2(new_n286), .A3(new_n324), .A4(new_n287), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n339), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n339), .A2(new_n345), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n288), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT79), .B1(new_n350), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n346), .A2(new_n286), .A3(new_n287), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n348), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n356), .A4(new_n355), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n288), .A2(new_n353), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n359), .ZN(new_n366));
  INV_X1    g165(.A(new_n356), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(new_n347), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n359), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n364), .A3(new_n356), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT82), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n370), .A3(new_n348), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n373), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n380), .A2(new_n381), .A3(new_n376), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n369), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G1gat), .B(G29gat), .Z(new_n384));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT6), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n388), .B(new_n369), .C1(new_n378), .C2(new_n382), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n375), .A2(KEYINPUT82), .A3(new_n377), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n381), .B1(new_n380), .B2(new_n376), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n396), .A2(KEYINPUT83), .A3(new_n388), .A4(new_n369), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n388), .B1(new_n396), .B2(new_n369), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G78gat), .B(G106gat), .Z(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT85), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406));
  NOR2_X1   g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407));
  AND2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408));
  AND2_X1   g207(.A1(G211gat), .A2(G218gat), .ZN(new_n409));
  OAI22_X1  g208(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(KEYINPUT22), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411));
  XOR2_X1   g210(.A(G211gat), .B(G218gat), .Z(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n410), .B(new_n412), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n406), .B(new_n413), .C1(new_n414), .C2(new_n411), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n346), .B1(new_n415), .B2(new_n351), .ZN(new_n416));
  AND2_X1   g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n406), .B2(new_n352), .ZN(new_n418));
  OR3_X1    g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n406), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n346), .B1(new_n420), .B2(new_n351), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n417), .B1(new_n421), .B2(new_n418), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT31), .B(G50gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n419), .B2(new_n422), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n405), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n404), .A3(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n227), .A2(new_n432), .A3(new_n277), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(KEYINPUT29), .ZN(new_n435));
  AOI211_X1 g234(.A(new_n414), .B(new_n434), .C1(new_n252), .C2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n414), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n280), .A2(new_n432), .A3(new_n228), .A4(new_n230), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n227), .A2(new_n277), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT74), .ZN(new_n443));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND4_X1  g245(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT30), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n438), .A2(new_n440), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n414), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n252), .A2(new_n435), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n437), .A3(new_n433), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT30), .A4(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n451), .ZN(new_n454));
  INV_X1    g253(.A(new_n446), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n447), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n454), .B2(new_n455), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n442), .A2(KEYINPUT75), .A3(new_n446), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n323), .A2(new_n401), .A3(new_n431), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n316), .A2(new_n321), .A3(new_n431), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n467), .A2(new_n466), .A3(new_n463), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n390), .A2(new_n393), .A3(new_n470), .A4(new_n397), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n400), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n465), .A2(new_n466), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n322), .A2(KEYINPUT36), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n316), .A2(new_n321), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n471), .A2(new_n400), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n463), .B1(new_n478), .B2(new_n469), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(new_n431), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n379), .A2(new_n355), .A3(new_n373), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n482), .A2(KEYINPUT87), .A3(new_n367), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT87), .B1(new_n482), .B2(new_n367), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n367), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(KEYINPUT87), .A3(new_n367), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n366), .A2(new_n367), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(new_n481), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n492), .A3(new_n388), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT40), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT88), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n399), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n463), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n493), .B2(KEYINPUT88), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n431), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n459), .A2(new_n460), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n446), .B1(new_n442), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n448), .B2(new_n437), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n450), .A2(new_n414), .A3(new_n433), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT38), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n398), .A2(KEYINPUT89), .A3(new_n400), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT38), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n454), .A2(KEYINPUT37), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n398), .A2(new_n400), .A3(new_n506), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n499), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n473), .B1(new_n480), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(G1gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT16), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519));
  OAI221_X1 g318(.A(new_n518), .B1(new_n519), .B2(G8gat), .C1(new_n517), .C2(new_n516), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(G8gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  XOR2_X1   g322(.A(G43gat), .B(G50gat), .Z(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n525), .A2(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n524), .B1(new_n530), .B2(KEYINPUT15), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(KEYINPUT15), .B2(new_n530), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n524), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n522), .B1(new_n523), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n533), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n535), .A2(new_n536), .B1(new_n534), .B2(new_n522), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n538), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n522), .B(new_n534), .Z(new_n543));
  XOR2_X1   g342(.A(new_n538), .B(KEYINPUT13), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G169gat), .B(G197gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n541), .A2(new_n542), .A3(new_n546), .A4(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT97), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT7), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n559), .A2(new_n561), .A3(G85gat), .A4(G92gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT97), .B(new_n558), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n562), .A2(new_n569), .A3(new_n565), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G57gat), .B(G64gat), .Z(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  INV_X1    g374(.A(G71gat), .ZN(new_n576));
  INV_X1    g375(.A(G78gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n574), .A2(new_n580), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n571), .A2(new_n582), .A3(new_n583), .A4(new_n572), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT98), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n588), .A3(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT100), .Z(new_n595));
  AND3_X1   g394(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n593), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT99), .B1(new_n590), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n591), .B(KEYINPUT101), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  NOR2_X1   g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  AOI211_X1 g405(.A(new_n592), .B(new_n606), .C1(new_n598), .C2(new_n591), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n522), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n584), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n584), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n611), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT20), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT93), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n616), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n534), .A2(new_n523), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n536), .A3(new_n573), .ZN(new_n628));
  INV_X1    g427(.A(new_n573), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT96), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n534), .A2(new_n629), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G190gat), .B(G218gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n608), .A2(new_n626), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n515), .A2(new_n557), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT102), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n515), .A2(new_n648), .A3(new_n557), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n469), .A2(new_n400), .A3(new_n471), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(KEYINPUT103), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(KEYINPUT103), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(G8gat), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT16), .B(G8gat), .Z(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n464), .B1(new_n647), .B2(new_n649), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n663), .B2(KEYINPUT105), .ZN(new_n664));
  INV_X1    g463(.A(new_n557), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n513), .A2(new_n507), .ZN(new_n666));
  INV_X1    g465(.A(new_n499), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n474), .A2(new_n476), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n472), .A2(new_n464), .ZN(new_n670));
  INV_X1    g469(.A(new_n431), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n665), .B1(new_n673), .B2(new_n473), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n648), .B1(new_n674), .B2(new_n645), .ZN(new_n675));
  INV_X1    g474(.A(new_n649), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n463), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n659), .B1(new_n664), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n663), .A2(KEYINPUT42), .A3(new_n661), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n657), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n659), .ZN(new_n684));
  OAI211_X1 g483(.A(KEYINPUT105), .B(new_n463), .C1(new_n675), .C2(new_n676), .ZN(new_n685));
  INV_X1    g484(.A(new_n662), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n663), .A2(KEYINPUT105), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(KEYINPUT106), .A3(new_n681), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n683), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n650), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n692), .A2(G15gat), .A3(new_n322), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n692), .B2(new_n477), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1326gat));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n692), .B2(new_n431), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n650), .A2(KEYINPUT107), .A3(new_n671), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n643), .ZN(new_n702));
  AND4_X1   g501(.A1(new_n674), .A2(new_n625), .A3(new_n702), .A4(new_n608), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n525), .A3(new_n654), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n643), .B1(new_n673), .B2(new_n473), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n515), .A2(new_n702), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n607), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n601), .B2(new_n604), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n665), .A2(new_n713), .A3(new_n626), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n652), .A2(new_n653), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n705), .A2(new_n717), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n528), .A3(new_n463), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT46), .Z(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n715), .B2(new_n464), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n711), .A2(new_n669), .A3(new_n714), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n322), .A2(G43gat), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n723), .A2(G43gat), .B1(new_n703), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g525(.A1(new_n703), .A2(new_n671), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n671), .A2(G50gat), .ZN(new_n728));
  OAI22_X1  g527(.A1(G50gat), .A2(new_n727), .B1(new_n715), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g529(.A1(new_n665), .A2(new_n626), .A3(new_n643), .A4(new_n713), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n673), .B2(new_n473), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n654), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g533(.A(new_n464), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT108), .Z(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n732), .A2(new_n576), .A3(new_n323), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n732), .A2(new_n669), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n576), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n671), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n557), .A2(new_n626), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n608), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n711), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n716), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n708), .B2(new_n747), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n746), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n654), .A2(new_n563), .A3(new_n713), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n755), .B2(new_n756), .ZN(G1336gat));
  NAND4_X1  g556(.A1(new_n707), .A2(new_n710), .A3(new_n463), .A4(new_n748), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n464), .A2(new_n608), .A3(G92gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n752), .A2(new_n753), .A3(new_n765), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT109), .B(new_n751), .C1(new_n708), .C2(new_n747), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n760), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n759), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(KEYINPUT52), .ZN(new_n770));
  AOI211_X1 g569(.A(KEYINPUT110), .B(new_n762), .C1(new_n768), .C2(new_n759), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n763), .B1(new_n770), .B2(new_n771), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n749), .B2(new_n477), .ZN(new_n773));
  OR3_X1    g572(.A1(new_n322), .A2(G99gat), .A3(new_n608), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n755), .B2(new_n774), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n608), .A2(G106gat), .A3(new_n431), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n766), .A2(new_n767), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n707), .A2(new_n710), .A3(new_n671), .A4(new_n748), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(G106gat), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT53), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  INV_X1    g580(.A(new_n776), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n755), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(new_n779), .ZN(G1339gat));
  OAI211_X1 g583(.A(new_n595), .B(new_n599), .C1(new_n596), .C2(new_n597), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n594), .B(KEYINPUT100), .ZN(new_n786));
  INV_X1    g585(.A(new_n597), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n593), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n591), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n785), .B(KEYINPUT54), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n598), .A2(new_n792), .A3(new_n600), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(new_n606), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n607), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n606), .A4(new_n793), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n702), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n547), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n537), .A2(new_n800), .A3(new_n538), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n537), .B2(new_n538), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n543), .A2(new_n803), .A3(new_n545), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n543), .A2(new_n545), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n801), .A2(new_n802), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n799), .A2(new_n553), .B1(new_n807), .B2(new_n552), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n798), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n811), .A2(new_n557), .A3(new_n712), .A4(new_n797), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n713), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n702), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n625), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n644), .A2(new_n557), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n716), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AND4_X1   g618(.A1(new_n431), .A2(new_n819), .A3(new_n464), .A4(new_n323), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n260), .A3(new_n557), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n671), .B1(new_n818), .B2(new_n815), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n323), .B1(new_n822), .B2(KEYINPUT114), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n716), .A2(new_n463), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n825), .A2(new_n557), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n821), .B1(new_n827), .B2(new_n260), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n821), .C1(new_n827), .C2(new_n260), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1340gat));
  NAND3_X1  g631(.A1(new_n820), .A2(new_n257), .A3(new_n713), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n825), .A2(new_n713), .A3(new_n826), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(G120gat), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n834), .B2(G120gat), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(G1341gat));
  NAND2_X1  g637(.A1(new_n825), .A2(new_n826), .ZN(new_n839));
  OAI21_X1  g638(.A(G127gat), .B1(new_n839), .B2(new_n625), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n253), .A3(new_n626), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  NAND4_X1  g641(.A1(new_n820), .A2(new_n265), .A3(new_n266), .A4(new_n702), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n839), .B2(new_n643), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n818), .A2(new_n815), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n848), .B2(new_n671), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n850), .B(new_n431), .C1(new_n818), .C2(new_n815), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n716), .A2(new_n463), .A3(new_n669), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G141gat), .B1(new_n854), .B2(new_n665), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n669), .A2(new_n431), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n665), .A2(G141gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n819), .A2(new_n464), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n819), .A2(new_n856), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(new_n463), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n857), .ZN(new_n865));
  XOR2_X1   g664(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n866));
  NAND2_X1  g665(.A1(new_n855), .A2(new_n866), .ZN(new_n867));
  OAI22_X1  g666(.A1(new_n859), .A2(new_n860), .B1(new_n865), .B2(new_n867), .ZN(G1344gat));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n869), .B(G148gat), .C1(new_n854), .C2(new_n608), .ZN(new_n870));
  INV_X1    g669(.A(new_n816), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n796), .A2(new_n872), .A3(new_n702), .A4(new_n797), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n808), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n798), .A2(KEYINPUT119), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n814), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(new_n626), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n877), .B2(new_n671), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n713), .B(new_n853), .C1(new_n878), .C2(new_n851), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G148gat), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n880), .B2(KEYINPUT59), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  AOI211_X1 g681(.A(new_n882), .B(new_n869), .C1(new_n879), .C2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n870), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n327), .A3(new_n713), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1345gat));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n331), .A3(new_n626), .ZN(new_n887));
  OAI21_X1  g686(.A(G155gat), .B1(new_n854), .B2(new_n625), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1346gat));
  NAND3_X1  g688(.A1(new_n864), .A2(new_n332), .A3(new_n702), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT121), .B1(new_n854), .B2(new_n643), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G162gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n854), .A2(KEYINPUT121), .A3(new_n643), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(G1347gat));
  AOI21_X1  g693(.A(new_n654), .B1(new_n815), .B2(new_n818), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n467), .A2(new_n464), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT122), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n557), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n654), .A2(new_n464), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n823), .A2(new_n824), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n665), .A2(new_n203), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n899), .A2(new_n901), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n713), .A2(new_n204), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n204), .B1(new_n906), .B2(new_n713), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT123), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n825), .A2(new_n904), .ZN(new_n914));
  OAI21_X1  g713(.A(G176gat), .B1(new_n914), .B2(new_n608), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n915), .B(new_n916), .C1(new_n909), .C2(new_n910), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n906), .A2(new_n626), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n626), .A2(new_n247), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n919), .A2(G183gat), .B1(new_n898), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  MUX2_X1   g722(.A(new_n923), .B(KEYINPUT60), .S(KEYINPUT125), .Z(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n921), .B2(new_n923), .ZN(G1350gat));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(G190gat), .C1(new_n914), .C2(new_n643), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n823), .A2(new_n824), .A3(new_n905), .A4(new_n643), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT126), .B1(new_n929), .B2(new_n223), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n930), .A3(KEYINPUT61), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  OAI211_X1 g731(.A(KEYINPUT126), .B(new_n932), .C1(new_n929), .C2(new_n223), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n902), .A2(new_n223), .A3(new_n702), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(G1351gat));
  AND3_X1   g734(.A1(new_n895), .A2(new_n463), .A3(new_n856), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n557), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n878), .A2(new_n851), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n904), .A2(new_n477), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n557), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n936), .A2(new_n943), .A3(new_n713), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT62), .Z(new_n945));
  NOR3_X1   g744(.A1(new_n938), .A2(new_n608), .A3(new_n939), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n943), .ZN(G1353gat));
  INV_X1    g746(.A(G211gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n936), .A2(new_n948), .A3(new_n626), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n940), .A2(new_n626), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  AOI21_X1  g752(.A(G218gat), .B1(new_n936), .B2(new_n702), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n702), .A2(G218gat), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT127), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n940), .B2(new_n956), .ZN(G1355gat));
endmodule


