//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT64), .A2(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n195), .A2(new_n191), .A3(new_n192), .A4(G214), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n190), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(KEYINPUT87), .A3(G131), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n201), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT86), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(new_n207), .A3(new_n201), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT88), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  XNOR2_X1  g026(.A(G125), .B(G140), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(KEYINPUT16), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT19), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n213), .B(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n219), .B2(KEYINPUT19), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n204), .A2(new_n223), .A3(new_n206), .A4(new_n208), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n210), .A2(new_n215), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT85), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n221), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n219), .A2(new_n229), .A3(G146), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n200), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n198), .A2(KEYINPUT18), .A3(G131), .A4(new_n199), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .A4(new_n205), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n189), .B1(new_n225), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n214), .B(new_n221), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n202), .A2(KEYINPUT17), .A3(new_n203), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n238), .B(new_n239), .C1(new_n209), .C2(KEYINPUT17), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n235), .A2(new_n189), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n244));
  INV_X1    g058(.A(G475), .ZN(new_n245));
  INV_X1    g059(.A(G902), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n245), .B(new_n246), .C1(new_n236), .C2(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT20), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n189), .B1(new_n235), .B2(new_n240), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n246), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G475), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT91), .A2(G952), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT91), .A2(G952), .ZN(new_n257));
  AOI21_X1  g071(.A(G953), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G234), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n191), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT21), .B(G898), .Z(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n246), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT9), .B(G234), .Z(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(G217), .A3(new_n192), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n268));
  INV_X1    g082(.A(G107), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT78), .A2(G107), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G116), .B(G122), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n196), .B2(new_n197), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(KEYINPUT67), .A2(G128), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT67), .A2(G128), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G143), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n277), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT13), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n277), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT89), .B1(new_n276), .B2(KEYINPUT13), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n281), .A4(new_n289), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n274), .B(new_n284), .C1(new_n290), .C2(G134), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n272), .A2(new_n273), .ZN(new_n292));
  INV_X1    g106(.A(G116), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT14), .A3(G122), .ZN(new_n294));
  INV_X1    g108(.A(new_n273), .ZN(new_n295));
  OAI211_X1 g109(.A(G107), .B(new_n294), .C1(new_n295), .C2(KEYINPUT14), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n282), .B1(new_n277), .B2(new_n281), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n292), .B(new_n296), .C1(new_n284), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n267), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n274), .B1(new_n290), .B2(G134), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n283), .ZN(new_n302));
  INV_X1    g116(.A(new_n267), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n304), .A3(KEYINPUT90), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT90), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n267), .C1(new_n291), .C2(new_n299), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n246), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G478), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n254), .A2(new_n265), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G221), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n266), .B2(new_n246), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n270), .A2(new_n188), .A3(new_n271), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT80), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n269), .A2(G104), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n270), .A2(new_n318), .A3(new_n188), .A4(new_n271), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT81), .ZN(new_n322));
  AND2_X1   g136(.A1(KEYINPUT64), .A2(G143), .ZN(new_n323));
  NOR2_X1   g137(.A1(KEYINPUT64), .A2(G143), .ZN(new_n324));
  OAI21_X1  g138(.A(G146), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n195), .A2(G146), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n325), .A2(new_n326), .A3(G128), .A4(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n196), .A2(new_n221), .A3(new_n197), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n275), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n196), .A2(new_n197), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(G146), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n272), .A2(new_n335), .A3(G104), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n269), .A2(G104), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(KEYINPUT3), .B2(new_n317), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n320), .A2(new_n341), .A3(G101), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n322), .A2(new_n334), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n320), .A2(new_n341), .A3(G101), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n320), .B2(G101), .ZN(new_n345));
  INV_X1    g159(.A(new_n340), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n221), .B2(G143), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n330), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n278), .B(new_n279), .C1(new_n327), .C2(new_n326), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n329), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n343), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT66), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G137), .ZN(new_n357));
  INV_X1    g171(.A(G137), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(KEYINPUT66), .ZN(new_n359));
  OAI211_X1 g173(.A(KEYINPUT11), .B(G134), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT11), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n282), .B2(G137), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n282), .A2(G137), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n360), .A2(new_n364), .A3(new_n201), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n201), .B1(new_n360), .B2(new_n364), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n355), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT12), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n325), .A2(G128), .A3(new_n328), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n371), .A2(new_n326), .B1(new_n351), .B2(new_n352), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n347), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n343), .A2(new_n373), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n336), .A2(new_n339), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT79), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n336), .A2(new_n380), .A3(new_n339), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n378), .A2(new_n379), .A3(G101), .A4(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT0), .B(G128), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n351), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n325), .A2(KEYINPUT0), .A3(G128), .A4(new_n328), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n336), .A2(new_n380), .A3(new_n339), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n380), .B1(new_n336), .B2(new_n339), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(new_n337), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n382), .B(new_n387), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n375), .A2(new_n376), .A3(new_n367), .A4(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G140), .ZN(new_n394));
  INV_X1    g208(.A(G227), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G953), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n394), .B(new_n396), .Z(new_n397));
  INV_X1    g211(.A(KEYINPUT12), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n355), .A2(new_n398), .A3(new_n368), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n370), .A2(new_n393), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT82), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n322), .A2(new_n340), .A3(new_n342), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n372), .ZN(new_n403));
  AOI211_X1 g217(.A(KEYINPUT12), .B(new_n367), .C1(new_n403), .C2(new_n343), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n398), .B1(new_n355), .B2(new_n368), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n393), .A4(new_n397), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n375), .A2(new_n376), .A3(new_n392), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n368), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n393), .ZN(new_n411));
  INV_X1    g225(.A(new_n397), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G469), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n246), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n246), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n410), .A2(new_n393), .A3(new_n397), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n370), .A2(new_n393), .A3(new_n399), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(G469), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n314), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G214), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT69), .B1(new_n293), .B2(G119), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT69), .ZN(new_n426));
  INV_X1    g240(.A(G119), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(G116), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n428), .C1(G116), .C2(new_n427), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT2), .B(G113), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n382), .B(new_n431), .C1(new_n390), .C2(new_n391), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n427), .A3(G116), .ZN(new_n434));
  OAI211_X1 g248(.A(G113), .B(new_n434), .C1(new_n429), .C2(new_n433), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n429), .A2(new_n430), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n322), .A2(new_n437), .A3(new_n340), .A4(new_n342), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(G110), .B(G122), .Z(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n440), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n442), .A3(new_n438), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n354), .A2(G125), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(G125), .B2(new_n386), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n192), .A2(G224), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n439), .A2(new_n449), .A3(new_n440), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(KEYINPUT7), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n446), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n402), .B(new_n437), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n440), .B(KEYINPUT8), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n443), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n246), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n451), .A2(new_n456), .A3(new_n246), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n424), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n312), .A2(new_n422), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n215), .A2(new_n228), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n275), .A2(G119), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n467), .A2(KEYINPUT75), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n280), .A2(G119), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT75), .ZN(new_n470));
  INV_X1    g284(.A(new_n467), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT24), .B(G110), .Z(new_n473));
  OR2_X1    g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n475), .B1(new_n427), .B2(G128), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n471), .B(new_n476), .C1(new_n469), .C2(new_n475), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n477), .A2(G110), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n466), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT22), .B(G137), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n313), .A2(new_n259), .A3(G953), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n238), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n472), .A2(new_n473), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n477), .A2(G110), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n483), .B(KEYINPUT76), .ZN(new_n489));
  INV_X1    g303(.A(new_n487), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n479), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n465), .B1(new_n492), .B2(new_n246), .ZN(new_n493));
  AOI211_X1 g307(.A(KEYINPUT25), .B(G902), .C1(new_n488), .C2(new_n491), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G217), .B1(new_n259), .B2(G902), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n496), .B(KEYINPUT74), .Z(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(G902), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT73), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n384), .B(new_n385), .C1(new_n365), .C2(new_n366), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n358), .A2(KEYINPUT66), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n356), .A2(G137), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n282), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n358), .A2(G134), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n201), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n362), .A2(new_n363), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n282), .B1(new_n504), .B2(new_n505), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(KEYINPUT11), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n508), .B1(new_n511), .B2(new_n201), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n354), .ZN(new_n513));
  INV_X1    g327(.A(new_n431), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n503), .A2(new_n513), .A3(new_n519), .A4(new_n514), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n503), .A2(new_n513), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n518), .A2(new_n520), .B1(new_n431), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n517), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n191), .A2(new_n192), .A3(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(G101), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n527), .B(KEYINPUT71), .Z(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(KEYINPUT68), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(KEYINPUT68), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n531), .B(new_n533), .C1(new_n503), .C2(new_n513), .ZN(new_n534));
  AND4_X1   g348(.A1(KEYINPUT68), .A2(new_n503), .A3(new_n513), .A4(new_n530), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n431), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n518), .A2(new_n520), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n527), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT31), .ZN(new_n539));
  INV_X1    g353(.A(new_n531), .ZN(new_n540));
  INV_X1    g354(.A(new_n366), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n360), .A2(new_n364), .A3(new_n201), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n386), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n506), .A2(new_n507), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G131), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n372), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n540), .B(new_n532), .C1(new_n543), .C2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n503), .A2(new_n513), .A3(KEYINPUT68), .A4(new_n530), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n550), .A2(new_n431), .B1(new_n518), .B2(new_n520), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT31), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n527), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n529), .A2(new_n539), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G472), .A2(G902), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n502), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(KEYINPUT73), .B(new_n557), .C1(new_n554), .C2(new_n555), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n551), .B2(new_n527), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n527), .B(new_n517), .C1(new_n522), .C2(new_n516), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n528), .A2(KEYINPUT29), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n523), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n246), .ZN(new_n569));
  INV_X1    g383(.A(new_n555), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n552), .B1(new_n551), .B2(new_n527), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n552), .A2(new_n536), .A3(new_n537), .A4(new_n527), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n573), .B2(new_n529), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n569), .A2(G472), .B1(new_n574), .B2(KEYINPUT32), .ZN(new_n575));
  AOI211_X1 g389(.A(KEYINPUT77), .B(new_n501), .C1(new_n561), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT73), .B1(new_n574), .B2(new_n557), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(G472), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(KEYINPUT32), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n556), .A2(new_n502), .A3(new_n558), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n501), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n464), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  NAND2_X1  g400(.A1(new_n416), .A2(new_n421), .ZN(new_n587));
  INV_X1    g401(.A(new_n314), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n501), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n554), .A2(new_n246), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT93), .Z(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n308), .A2(new_n309), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n308), .A2(KEYINPUT94), .A3(new_n309), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n305), .A2(new_n603), .A3(new_n307), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n300), .A2(new_n304), .A3(KEYINPUT33), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n309), .A2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n254), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n457), .A2(new_n458), .ZN(new_n611));
  INV_X1    g425(.A(new_n265), .ZN(new_n612));
  INV_X1    g426(.A(new_n458), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n451), .A2(new_n456), .A3(new_n246), .A4(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n611), .A2(new_n423), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n597), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n188), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  NAND2_X1  g434(.A1(new_n311), .A2(new_n253), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n622));
  OR3_X1    g436(.A1(new_n248), .A2(new_n622), .A3(KEYINPUT20), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n622), .B1(new_n248), .B2(KEYINPUT20), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n249), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(KEYINPUT97), .A3(new_n249), .A4(new_n624), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n621), .B(new_n615), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n597), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND2_X1  g446(.A1(new_n480), .A2(new_n487), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT98), .ZN(new_n634));
  INV_X1    g448(.A(new_n489), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n636));
  OR3_X1    g450(.A1(new_n479), .A2(new_n490), .A3(KEYINPUT98), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n499), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n498), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n464), .A2(new_n594), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G110), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  AND3_X1   g460(.A1(new_n611), .A2(new_n423), .A3(new_n614), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n642), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n582), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n628), .ZN(new_n650));
  INV_X1    g464(.A(new_n264), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT100), .B(G900), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n260), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT101), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n621), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n650), .A2(new_n422), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n275), .ZN(G30));
  INV_X1    g472(.A(new_n522), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n528), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n538), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n246), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n660), .B2(new_n538), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n578), .A2(new_n580), .A3(new_n581), .A4(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n561), .A2(KEYINPUT103), .A3(new_n580), .A4(new_n665), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n642), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n654), .B(KEYINPUT39), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n422), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT104), .Z(new_n674));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n673), .B(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n460), .A2(new_n462), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT38), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n247), .A2(new_n249), .B1(G475), .B2(new_n252), .ZN(new_n681));
  INV_X1    g495(.A(new_n311), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n680), .A2(new_n423), .A3(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n670), .A2(new_n676), .A3(new_n678), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n332), .ZN(G45));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n600), .A2(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n681), .A2(new_n688), .A3(new_n654), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n422), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n687), .B1(new_n649), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n690), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n647), .A2(new_n642), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n561), .B2(new_n575), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n694), .A3(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  AOI21_X1  g511(.A(new_n501), .B1(new_n561), .B2(new_n575), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n414), .A2(new_n415), .A3(new_n246), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n415), .B1(new_n414), .B2(new_n246), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n699), .B1(new_n702), .B2(new_n588), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT106), .A4(new_n314), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n698), .B(new_n616), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  OAI211_X1 g521(.A(new_n698), .B(new_n629), .C1(new_n703), .C2(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR3_X1   g523(.A1(new_n700), .A2(new_n701), .A3(new_n314), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n694), .A2(new_n312), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT107), .B(G119), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G21));
  NAND3_X1  g527(.A1(new_n683), .A2(new_n647), .A3(new_n612), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n591), .A2(G472), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n583), .A2(new_n556), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n703), .B2(new_n704), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  AND3_X1   g533(.A1(new_n642), .A2(new_n715), .A3(new_n556), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n710), .A2(new_n647), .A3(new_n689), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  NAND3_X1  g536(.A1(new_n460), .A2(new_n423), .A3(new_n462), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n574), .A2(KEYINPUT32), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n501), .B1(new_n575), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n582), .A2(new_n583), .A3(new_n724), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(new_n690), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n692), .A2(new_n698), .A3(KEYINPUT108), .A4(new_n724), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n727), .B1(new_n732), .B2(KEYINPUT42), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  AND3_X1   g548(.A1(new_n650), .A2(new_n422), .A3(new_n655), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n698), .A3(new_n724), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n609), .A2(new_n681), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT43), .ZN(new_n739));
  INV_X1    g553(.A(new_n642), .ZN(new_n740));
  OR3_X1    g554(.A1(new_n739), .A2(new_n594), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n723), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n420), .A2(KEYINPUT45), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n397), .B1(new_n406), .B2(new_n393), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n747), .B2(new_n418), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n748), .A3(G469), .ZN(new_n749));
  INV_X1    g563(.A(new_n417), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n416), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n588), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n671), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT109), .B1(new_n741), .B2(new_n742), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n741), .A2(KEYINPUT109), .A3(new_n742), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n744), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n588), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n582), .A2(new_n583), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n689), .A3(new_n724), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NOR2_X1   g582(.A1(new_n739), .A2(new_n260), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n700), .A2(new_n701), .A3(new_n723), .A4(new_n314), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n726), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT48), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n739), .A2(new_n260), .A3(new_n716), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n680), .A2(new_n423), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n710), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n501), .A2(new_n260), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n668), .A2(new_n669), .A3(new_n770), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n681), .A3(new_n688), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n773), .A2(new_n724), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n702), .A2(KEYINPUT114), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n702), .A2(KEYINPUT114), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n314), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT115), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(new_n314), .C1(new_n784), .C2(new_n785), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n783), .B1(new_n765), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n769), .A2(new_n720), .A3(new_n770), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT116), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n777), .A2(new_n782), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n773), .A2(new_n647), .A3(new_n710), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n779), .B(KEYINPUT117), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n258), .B(new_n797), .C1(new_n798), .C2(new_n610), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n781), .A2(new_n254), .A3(new_n609), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n258), .A4(new_n797), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n763), .A2(new_n764), .A3(new_n786), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n795), .B1(new_n805), .B2(new_n783), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n777), .A2(new_n806), .A3(new_n782), .A4(new_n793), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n772), .A2(new_n796), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n721), .B1(new_n649), .B2(new_n656), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n691), .B2(new_n695), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n668), .A2(new_n669), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n423), .A2(new_n683), .A3(new_n614), .A4(new_n611), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n589), .A2(new_n654), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n740), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n414), .A2(new_n246), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(G469), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n647), .A3(new_n588), .A4(new_n416), .ZN(new_n818));
  INV_X1    g632(.A(new_n654), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n254), .A2(new_n609), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n735), .A2(new_n694), .B1(new_n821), .B2(new_n720), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n696), .A2(new_n814), .A3(KEYINPUT52), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n815), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n610), .B1(new_n254), .B2(new_n682), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n463), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n612), .A3(new_n590), .A4(new_n594), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n585), .A2(new_n828), .A3(new_n708), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n643), .A2(new_n705), .A3(new_n711), .A4(new_n718), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n720), .A2(new_n422), .A3(new_n689), .A4(new_n724), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT111), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n682), .A2(new_n253), .A3(new_n819), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n582), .A2(new_n422), .A3(new_n650), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n724), .A2(new_n642), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n834), .A2(new_n835), .B1(new_n729), .B2(new_n656), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n733), .A2(new_n829), .A3(new_n830), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n825), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(KEYINPUT112), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n824), .A2(KEYINPUT113), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n696), .A2(new_n814), .A3(new_n822), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n823), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n838), .B2(KEYINPUT112), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT54), .B(new_n839), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n825), .B2(new_n838), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n733), .A2(new_n829), .A3(new_n830), .A4(new_n837), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n846), .A3(KEYINPUT53), .A4(new_n841), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n808), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(G952), .A2(G953), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n808), .A2(new_n850), .A3(KEYINPUT119), .A4(new_n855), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT49), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n583), .B(new_n588), .C1(new_n702), .C2(new_n862), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n863), .A2(new_n424), .A3(new_n738), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n680), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n811), .B1(new_n862), .B2(new_n702), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n861), .A2(new_n870), .ZN(G75));
  AOI21_X1  g685(.A(new_n246), .B1(new_n851), .B2(new_n853), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT56), .B1(new_n872), .B2(G210), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n444), .A2(new_n450), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n448), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT55), .Z(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n873), .A2(new_n877), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n192), .A2(G952), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G51));
  XNOR2_X1  g695(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n417), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n854), .B1(new_n851), .B2(new_n853), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT121), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n414), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n749), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n880), .B1(new_n890), .B2(new_n892), .ZN(G54));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n245), .A3(KEYINPUT122), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n246), .B(new_n895), .C1(new_n851), .C2(new_n853), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT122), .B1(new_n894), .B2(new_n245), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n243), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n899));
  INV_X1    g713(.A(new_n895), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n872), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n243), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n896), .A2(KEYINPUT123), .A3(new_n243), .A4(new_n897), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n880), .B(new_n898), .C1(new_n903), .C2(new_n904), .ZN(G60));
  XNOR2_X1  g719(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n309), .A2(new_n246), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n906), .B(new_n907), .Z(new_n908));
  OAI211_X1 g722(.A(new_n606), .B(new_n908), .C1(new_n884), .C2(new_n885), .ZN(new_n909));
  INV_X1    g723(.A(new_n880), .ZN(new_n910));
  INV_X1    g724(.A(new_n908), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n850), .B2(new_n855), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n909), .B(new_n910), .C1(new_n912), .C2(new_n606), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(new_n851), .A2(new_n853), .ZN(new_n915));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  NOR2_X1   g731(.A1(new_n639), .A2(new_n640), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT125), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n910), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n492), .B1(new_n915), .B2(new_n917), .ZN(new_n923));
  OR3_X1    g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  NAND2_X1  g740(.A1(new_n829), .A2(new_n830), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n192), .B1(new_n262), .B2(G224), .ZN(new_n929));
  AOI22_X1  g743(.A1(new_n927), .A2(new_n192), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n874), .B1(G898), .B2(new_n192), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  NAND3_X1  g747(.A1(new_n757), .A2(new_n726), .A3(new_n812), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n767), .A2(new_n810), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n733), .A2(new_n736), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n760), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT127), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n939), .A3(new_n760), .A4(new_n936), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n192), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n550), .B(new_n220), .ZN(new_n942));
  INV_X1    g756(.A(G900), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n943), .B2(G227), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n810), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n685), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n760), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n826), .A2(new_n724), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n674), .B(new_n951), .C1(new_n584), .C2(new_n576), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n767), .B(new_n952), .C1(new_n947), .C2(new_n948), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n192), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n942), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n395), .B2(new_n943), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n945), .A2(new_n957), .ZN(G72));
  INV_X1    g772(.A(new_n551), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(new_n527), .ZN(new_n960));
  INV_X1    g774(.A(new_n927), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n938), .A2(new_n961), .A3(new_n940), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n960), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n959), .A2(new_n527), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n950), .A2(new_n953), .A3(new_n927), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n965), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n910), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n839), .B1(new_n847), .B2(new_n849), .ZN(new_n971));
  NOR4_X1   g785(.A1(new_n971), .A2(new_n965), .A3(new_n967), .A4(new_n960), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(G57));
endmodule


