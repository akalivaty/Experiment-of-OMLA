//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G214), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT18), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n193), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G237), .ZN(new_n200));
  INV_X1    g014(.A(G953), .ZN(new_n201));
  AND4_X1   g015(.A1(G143), .A2(new_n200), .A3(new_n201), .A4(G214), .ZN(new_n202));
  AOI21_X1  g016(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n204), .B(KEYINPUT92), .C1(new_n195), .C2(new_n196), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT73), .B1(new_n208), .B2(G140), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(KEYINPUT74), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n217), .A3(G140), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n207), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(G125), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n208), .A2(G140), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n207), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT91), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n218), .ZN(new_n225));
  OAI21_X1  g039(.A(G146), .B1(new_n225), .B2(new_n213), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n222), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n202), .B2(new_n203), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT18), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n206), .A2(new_n224), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n218), .A2(KEYINPUT16), .A3(new_n209), .A4(new_n212), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n215), .A2(new_n217), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT16), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n211), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(G146), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(G146), .B1(new_n233), .B2(new_n236), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI211_X1 g055(.A(new_n238), .B(G146), .C1(new_n233), .C2(new_n236), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT95), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n204), .A2(new_n196), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n229), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n246), .B2(KEYINPUT17), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n245), .A2(KEYINPUT95), .A3(new_n248), .A4(new_n229), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n189), .B(new_n232), .C1(new_n243), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n237), .A2(KEYINPUT77), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT19), .B1(new_n225), .B2(new_n213), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT19), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n220), .A2(new_n221), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT93), .ZN(new_n257));
  OR2_X1    g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n254), .A2(new_n258), .A3(new_n207), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n233), .A2(new_n261), .A3(new_n236), .A4(G146), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n253), .A2(new_n260), .A3(new_n262), .A4(new_n246), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT94), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n232), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n189), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n232), .B2(new_n263), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n252), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n270));
  NOR2_X1   g084(.A1(G475), .A2(G902), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT96), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT97), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT97), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n269), .A2(new_n276), .A3(new_n270), .A4(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n273), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT20), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n232), .B1(new_n243), .B2(new_n251), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n282), .A2(new_n266), .ZN(new_n283));
  INV_X1    g097(.A(new_n252), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G475), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n281), .B(new_n201), .C1(G234), .C2(G237), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT21), .B(G898), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(KEYINPUT101), .A2(G952), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT101), .A2(G952), .ZN(new_n292));
  AOI21_X1  g106(.A(G953), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G234), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n200), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G107), .ZN(new_n297));
  INV_X1    g111(.A(G116), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n298), .A2(G122), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(KEYINPUT14), .ZN(new_n300));
  XNOR2_X1  g114(.A(G116), .B(G122), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n300), .A2(new_n303), .B1(new_n297), .B2(new_n301), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT98), .ZN(new_n305));
  INV_X1    g119(.A(G128), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(G143), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n192), .A2(KEYINPUT98), .A3(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G134), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(G143), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(KEYINPUT99), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n301), .B(new_n297), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT99), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n309), .A2(new_n318), .A3(new_n310), .A4(new_n311), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT13), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n309), .A2(new_n321), .B1(new_n306), .B2(G143), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n307), .A2(KEYINPUT13), .A3(new_n308), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n310), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n315), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT9), .B(G234), .ZN(new_n326));
  INV_X1    g140(.A(G217), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(G953), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n315), .B(new_n328), .C1(new_n320), .C2(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT100), .B1(new_n332), .B2(new_n281), .ZN(new_n333));
  INV_X1    g147(.A(G478), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(KEYINPUT15), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT100), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n337), .B(G902), .C1(new_n330), .C2(new_n331), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n287), .A2(new_n296), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G214), .B1(G237), .B2(G902), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT88), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n188), .A2(KEYINPUT3), .A3(G107), .ZN(new_n344));
  AND2_X1   g158(.A1(KEYINPUT83), .A2(G104), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT83), .A2(G104), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n297), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT85), .B(G101), .Z(new_n349));
  NOR2_X1   g163(.A1(new_n345), .A2(new_n346), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT84), .B1(new_n350), .B2(G107), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n352));
  NOR4_X1   g166(.A1(new_n345), .A2(new_n346), .A3(new_n352), .A4(new_n297), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n348), .B(new_n349), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT4), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  OR2_X1    g170(.A1(KEYINPUT83), .A2(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT83), .A2(G104), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(G107), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n352), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n350), .A2(KEYINPUT84), .A3(G107), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(new_n362), .B2(new_n348), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT86), .B1(new_n355), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G101), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT4), .A4(new_n354), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  OR3_X1    g183(.A1(new_n298), .A2(KEYINPUT66), .A3(G119), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT66), .B1(new_n298), .B2(G119), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n298), .A2(G119), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT2), .B(G113), .Z(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n376), .A3(G101), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n363), .A2(KEYINPUT87), .A3(new_n376), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n369), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n347), .B1(G104), .B2(new_n297), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n354), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n373), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT5), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n298), .A2(KEYINPUT5), .A3(G119), .ZN(new_n389));
  INV_X1    g203(.A(G113), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n388), .A2(new_n391), .B1(new_n374), .B2(new_n387), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G122), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT89), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT0), .A2(G128), .ZN(new_n402));
  XNOR2_X1  g216(.A(G143), .B(G146), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n207), .A2(G143), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n192), .A2(G146), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT0), .B(G128), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT64), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n234), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n413));
  OAI21_X1  g227(.A(G128), .B1(new_n413), .B2(KEYINPUT65), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n406), .B2(KEYINPUT1), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n408), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n403), .A2(new_n418), .A3(G128), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n412), .B1(new_n421), .B2(new_n234), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n201), .A2(G224), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n382), .A2(new_n394), .A3(new_n397), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT6), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n399), .B1(new_n382), .B2(new_n394), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n401), .B(new_n424), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(KEYINPUT7), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n412), .B(new_n429), .C1(new_n421), .C2(new_n234), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT90), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n422), .A2(KEYINPUT7), .A3(new_n423), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n397), .B(KEYINPUT8), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n386), .A2(new_n392), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n393), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n436), .B2(new_n425), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n437), .A3(new_n439), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n343), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G221), .B1(new_n326), .B2(G902), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT81), .Z(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n281), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n306), .B1(new_n406), .B2(KEYINPUT1), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n419), .B1(new_n448), .B2(new_n403), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n354), .A2(new_n384), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n354), .A2(new_n420), .A3(KEYINPUT10), .A4(new_n384), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n411), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n379), .B2(new_n380), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n369), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n310), .B2(G137), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n310), .A2(G137), .ZN(new_n460));
  INV_X1    g274(.A(G137), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT11), .A3(G134), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G131), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n459), .A2(new_n462), .A3(new_n196), .A4(new_n460), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n457), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n385), .A2(new_n421), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n469), .B2(new_n450), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT12), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  INV_X1    g287(.A(G227), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n473), .B(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT82), .Z(new_n477));
  AND2_X1   g291(.A1(new_n369), .A2(new_n456), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n466), .B1(new_n478), .B2(new_n454), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n457), .B2(new_n467), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n472), .A2(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n447), .B1(new_n481), .B2(G469), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n457), .A2(new_n467), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n466), .B(new_n454), .C1(new_n369), .C2(new_n456), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n480), .A2(new_n471), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n446), .A3(new_n281), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n445), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n341), .A2(new_n443), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n306), .A2(G119), .ZN(new_n494));
  INV_X1    g308(.A(G119), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT24), .B(G110), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT76), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n306), .A2(KEYINPUT23), .A3(G119), .ZN(new_n503));
  INV_X1    g317(.A(G110), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n496), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT76), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n253), .A2(new_n262), .A3(new_n508), .A4(new_n222), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT78), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n508), .A2(new_n222), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(KEYINPUT78), .A3(new_n253), .A4(new_n262), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n241), .ZN(new_n515));
  INV_X1    g329(.A(new_n242), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n497), .A2(new_n498), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n502), .A2(new_n503), .A3(new_n496), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(G110), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n201), .A2(G221), .A3(G234), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n514), .B2(new_n520), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n493), .B1(new_n527), .B2(new_n281), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n514), .A2(new_n520), .ZN(new_n529));
  INV_X1    g343(.A(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n531), .A2(new_n493), .A3(new_n281), .A4(new_n524), .ZN(new_n532));
  OAI21_X1  g346(.A(G217), .B1(new_n294), .B2(G902), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT72), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n492), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n281), .A3(new_n524), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT25), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT79), .A3(new_n532), .A4(new_n535), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n527), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT80), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT80), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n537), .A2(new_n545), .A3(new_n542), .A4(new_n540), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT26), .B(G101), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n190), .A2(G210), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n553));
  NOR2_X1   g367(.A1(new_n461), .A2(G134), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n310), .A2(G137), .ZN(new_n555));
  OAI21_X1  g369(.A(G131), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n465), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n420), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n466), .A2(KEYINPUT67), .A3(new_n411), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT67), .B1(new_n466), .B2(new_n411), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n375), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n557), .B1(new_n417), .B2(new_n419), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n465), .A2(new_n464), .B1(new_n405), .B2(new_n410), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(new_n375), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n553), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n466), .A2(new_n411), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n375), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n552), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT30), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT67), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n466), .A2(new_n411), .A3(KEYINPUT67), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n564), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT30), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n563), .B1(new_n583), .B2(new_n572), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT31), .B1(new_n584), .B2(new_n552), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n576), .B1(new_n586), .B2(KEYINPUT30), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n552), .B(new_n562), .C1(new_n587), .C2(new_n375), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT31), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n575), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(G472), .A2(G902), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(KEYINPUT32), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT71), .ZN(new_n594));
  INV_X1    g408(.A(new_n592), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n583), .A2(new_n572), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(KEYINPUT31), .A3(new_n552), .A4(new_n562), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n595), .B1(new_n599), .B2(new_n575), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT71), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT32), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  INV_X1    g418(.A(new_n584), .ZN(new_n605));
  INV_X1    g419(.A(new_n552), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT29), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n568), .A2(new_n552), .A3(new_n573), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n586), .A2(new_n572), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n562), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT28), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n613), .A2(new_n573), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n606), .A2(new_n608), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n604), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n574), .B1(new_n596), .B2(new_n598), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n595), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT70), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(KEYINPUT70), .B(new_n619), .C1(new_n620), .C2(new_n595), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n603), .A2(new_n618), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n491), .A2(new_n547), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(new_n349), .Z(G3));
  NOR2_X1   g441(.A1(new_n332), .A2(KEYINPUT33), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n325), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n328), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n331), .A2(KEYINPUT104), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n325), .B(new_n629), .C1(KEYINPUT104), .C2(new_n329), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n628), .B1(new_n635), .B2(KEYINPUT33), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n334), .A2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n332), .A2(new_n281), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n637), .A2(new_n638), .B1(new_n334), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n280), .B2(new_n286), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n343), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n428), .A2(new_n437), .A3(new_n439), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n439), .B1(new_n428), .B2(new_n437), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT102), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n648), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n296), .B(new_n642), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n591), .A2(new_n281), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n600), .B1(new_n651), .B2(G472), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n544), .A2(new_n546), .A3(new_n489), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  AOI21_X1  g471(.A(new_n296), .B1(new_n647), .B2(new_n649), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n270), .B1(new_n269), .B2(new_n273), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n279), .A2(KEYINPUT105), .A3(new_n274), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n286), .A2(new_n662), .A3(new_n663), .A4(new_n340), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n654), .A2(new_n658), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NOR2_X1   g481(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n529), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n541), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n537), .A2(new_n540), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n652), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n490), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n647), .A2(new_n649), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n625), .ZN(new_n677));
  OR2_X1    g491(.A1(KEYINPUT106), .A2(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(KEYINPUT106), .A2(G900), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n288), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n295), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n489), .A2(new_n664), .A3(new_n671), .A4(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT107), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n601), .B1(new_n600), .B2(KEYINPUT32), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n620), .A2(KEYINPUT71), .A3(new_n619), .A4(new_n595), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n623), .B(new_n624), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n688), .A2(new_n618), .B1(new_n647), .B2(new_n649), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n682), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XNOR2_X1  g507(.A(new_n681), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n489), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT108), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n605), .A2(new_n552), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n612), .A2(new_n552), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(G902), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n604), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n687), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n441), .A2(new_n442), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT38), .ZN(new_n705));
  INV_X1    g519(.A(new_n671), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n287), .A2(new_n340), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n643), .A2(new_n705), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n697), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  NAND2_X1  g524(.A1(new_n489), .A2(new_n671), .ZN(new_n711));
  INV_X1    g525(.A(new_n640), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n287), .A2(new_n712), .A3(new_n681), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n689), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  OAI211_X1 g530(.A(new_n544), .B(new_n546), .C1(new_n687), .C2(new_n617), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n487), .A2(new_n281), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n444), .A3(new_n488), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n650), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT109), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n722), .B(new_n724), .ZN(G15));
  NAND4_X1  g539(.A1(new_n662), .A2(new_n663), .A3(new_n286), .A4(new_n340), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n296), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n544), .A2(new_n727), .A3(new_n546), .ZN(new_n728));
  INV_X1    g542(.A(new_n720), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n625), .A3(new_n676), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  AND2_X1   g545(.A1(new_n341), .A2(new_n671), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n676), .A3(new_n625), .A4(new_n729), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  NAND2_X1  g548(.A1(new_n651), .A2(G472), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n599), .B1(new_n552), .B2(new_n614), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n592), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n543), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n720), .A2(new_n296), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n676), .A2(new_n707), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  AOI21_X1  g556(.A(new_n720), .B1(new_n647), .B2(new_n649), .ZN(new_n743));
  INV_X1    g557(.A(new_n681), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n744), .B(new_n640), .C1(new_n286), .C2(new_n280), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n651), .A2(G472), .B1(new_n736), .B2(new_n592), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n671), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NOR3_X1   g564(.A1(new_n644), .A2(new_n645), .A3(new_n343), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n482), .A2(new_n488), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n444), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n717), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  AOI211_X1 g570(.A(G469), .B(G902), .C1(new_n485), .C2(new_n486), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT12), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n470), .B(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n477), .B1(new_n484), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n480), .A2(new_n479), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(G469), .ZN(new_n762));
  INV_X1    g576(.A(new_n447), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n444), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n441), .A2(new_n643), .A3(new_n442), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n765), .A2(new_n713), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n617), .B1(KEYINPUT32), .B2(new_n600), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n543), .B1(new_n768), .B2(new_n621), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n754), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n756), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  INV_X1    g586(.A(new_n717), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n726), .A2(new_n744), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n765), .A2(new_n766), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(KEYINPUT110), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n625), .A2(new_n775), .A3(new_n544), .A4(new_n546), .ZN(new_n778));
  INV_X1    g592(.A(new_n774), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  OAI21_X1  g596(.A(G469), .B1(new_n481), .B2(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(KEYINPUT45), .B2(new_n481), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n447), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n488), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n444), .B(new_n694), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n706), .A2(new_n652), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n287), .A2(new_n640), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT43), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT111), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(KEYINPUT111), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n788), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n751), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(KEYINPUT112), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(KEYINPUT112), .B2(new_n798), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT113), .B(G137), .Z(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(G39));
  OAI21_X1  g616(.A(new_n444), .B1(new_n786), .B2(new_n787), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT47), .Z(new_n804));
  NOR4_X1   g618(.A1(new_n547), .A2(new_n625), .A3(new_n713), .A4(new_n766), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  INV_X1    g621(.A(new_n295), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n791), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n739), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n743), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n720), .A2(new_n766), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n547), .A2(new_n808), .A3(new_n702), .A4(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(new_n642), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n293), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n811), .A2(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n769), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT48), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(new_n671), .A3(new_n746), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n815), .A2(new_n287), .A3(new_n712), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n719), .A2(new_n445), .A3(new_n488), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n751), .B(new_n812), .C1(new_n804), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(KEYINPUT121), .A2(KEYINPUT50), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n705), .A2(new_n643), .A3(new_n720), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n812), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n830), .B1(new_n812), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n822), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT122), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n812), .A2(new_n831), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n829), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n832), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n827), .B(new_n825), .C1(new_n838), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n836), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n676), .A2(new_n625), .A3(new_n729), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n846), .A2(new_n728), .B1(new_n721), .B2(new_n650), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n648), .B1(new_n704), .B2(new_n643), .ZN(new_n848));
  INV_X1    g662(.A(new_n649), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n707), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n740), .A2(new_n739), .ZN(new_n851));
  INV_X1    g665(.A(new_n296), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n340), .A2(KEYINPUT116), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n336), .A2(new_n339), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n287), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n443), .B(new_n852), .C1(new_n857), .C2(new_n641), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n850), .A2(new_n851), .B1(new_n653), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n490), .B1(new_n717), .B2(new_n672), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n847), .A2(new_n861), .A3(new_n733), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n681), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n662), .A2(new_n663), .A3(new_n286), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n751), .A3(new_n489), .A4(new_n671), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n687), .A2(new_n617), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n866), .A2(new_n867), .B1(new_n747), .B2(new_n753), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n756), .A2(new_n868), .A3(new_n770), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n781), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n845), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n689), .A2(new_n714), .B1(new_n743), .B2(new_n748), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n765), .A2(new_n671), .A3(new_n744), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n703), .A2(new_n676), .A3(new_n707), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n690), .B1(new_n689), .B2(new_n682), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n690), .A2(new_n682), .A3(new_n676), .A4(new_n625), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n872), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n692), .A2(KEYINPUT52), .A3(new_n872), .A4(new_n874), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n547), .A2(new_n625), .A3(new_n775), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n745), .A2(new_n751), .A3(new_n444), .A4(new_n752), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n618), .A2(new_n593), .A3(new_n621), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n537), .A3(new_n540), .A4(new_n542), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT42), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n748), .A2(new_n775), .ZN(new_n888));
  INV_X1    g702(.A(new_n711), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n625), .A3(new_n751), .A4(new_n865), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n883), .A2(new_n887), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n780), .B2(new_n776), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n658), .A2(new_n641), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n547), .A2(new_n625), .A3(new_n729), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n730), .B(new_n733), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n653), .A2(new_n858), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n626), .A3(new_n673), .A4(new_n741), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n898), .A3(KEYINPUT117), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n871), .A2(new_n881), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n881), .A2(KEYINPUT53), .A3(new_n898), .A4(new_n892), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n900), .A2(KEYINPUT119), .A3(new_n903), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT119), .B1(new_n900), .B2(new_n903), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n844), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(G952), .A2(G953), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n543), .A2(new_n343), .A3(new_n445), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n790), .B1(new_n914), .B2(KEYINPUT114), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(KEYINPUT114), .B2(new_n914), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n719), .A2(new_n488), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT49), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n703), .A2(new_n921), .A3(new_n705), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n913), .A2(new_n923), .ZN(G75));
  OAI21_X1  g738(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(G210), .A3(G902), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n401), .B1(new_n426), .B2(new_n427), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n424), .Z(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n926), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n926), .B2(new_n927), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n201), .A2(G952), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G51));
  XNOR2_X1  g750(.A(new_n447), .B(KEYINPUT57), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n900), .A2(new_n903), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n900), .A2(KEYINPUT119), .A3(new_n903), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n906), .B1(new_n942), .B2(new_n907), .ZN(new_n943));
  INV_X1    g757(.A(new_n910), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n487), .B(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n925), .A2(G902), .A3(new_n784), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n935), .B1(new_n947), .B2(new_n948), .ZN(G54));
  INV_X1    g763(.A(new_n935), .ZN(new_n950));
  AND2_X1   g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n925), .A2(G902), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(new_n269), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n925), .A2(G902), .A3(new_n269), .A4(new_n951), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(KEYINPUT125), .A3(new_n269), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G60));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n910), .B2(new_n905), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(new_n637), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n636), .A2(new_n960), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n910), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n962), .A2(new_n965), .A3(new_n935), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT126), .Z(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT60), .Z(new_n969));
  NAND3_X1  g783(.A1(new_n925), .A2(new_n669), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n942), .B2(new_n907), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n970), .B(new_n950), .C1(new_n972), .C2(new_n527), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n925), .A2(new_n969), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n525), .B2(new_n526), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n950), .A4(new_n970), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(new_n978), .ZN(G66));
  INV_X1    g793(.A(G224), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n289), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n898), .B2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n928), .B1(G898), .B2(new_n201), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G69));
  INV_X1    g798(.A(new_n806), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n642), .B1(new_n287), .B2(new_n856), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n773), .A2(new_n696), .A3(new_n751), .A4(new_n986), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n800), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n692), .A2(new_n872), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n709), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT62), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n254), .A2(new_n258), .A3(new_n259), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n583), .B(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n201), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(G900), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n994), .B2(new_n474), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n676), .A2(new_n707), .A3(new_n769), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n771), .B1(new_n788), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n985), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n781), .A3(new_n989), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n1001), .A2(G953), .A3(new_n800), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(G227), .B2(G953), .ZN(new_n1003));
  OAI221_X1 g817(.A(new_n995), .B1(new_n201), .B2(new_n997), .C1(new_n1003), .C2(new_n994), .ZN(G72));
  NAND3_X1  g818(.A1(new_n988), .A2(new_n898), .A3(new_n991), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  AOI21_X1  g821(.A(new_n698), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1000), .A2(new_n781), .A3(new_n989), .A4(new_n898), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1007), .B1(new_n1009), .B2(new_n800), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1010), .A2(new_n606), .A3(new_n584), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n607), .B(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n588), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n904), .A2(new_n1007), .A3(new_n1013), .ZN(new_n1014));
  NOR4_X1   g828(.A1(new_n1008), .A2(new_n1011), .A3(new_n935), .A4(new_n1014), .ZN(G57));
endmodule


