//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  OR2_X1    g0011(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n212), .A2(G50), .A3(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n220), .B1(new_n221), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n223), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n202), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT67), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n235));
  AOI22_X1  g0035(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n232), .A2(new_n233), .ZN(new_n238));
  OAI21_X1  g0038(.A(new_n221), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g0039(.A(new_n219), .B(new_n227), .C1(new_n239), .C2(KEYINPUT1), .ZN(new_n240));
  AOI21_X1  g0040(.A(new_n240), .B1(KEYINPUT1), .B2(new_n239), .ZN(G361));
  XOR2_X1   g0041(.A(G238), .B(G244), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XOR2_X1   g0047(.A(G264), .B(G270), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n245), .B(new_n249), .Z(G358));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT69), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G68), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G87), .B(G97), .Z(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(G200), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1698), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G222), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(G1698), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n265), .B1(new_n230), .B2(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n274), .A2(G274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n216), .ZN(new_n279));
  NAND3_X1  g0079(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n216), .B1(new_n277), .B2(new_n276), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n274), .B1(new_n284), .B2(new_n280), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(G226), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n259), .B1(new_n271), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n271), .A2(new_n286), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(G190), .ZN(new_n290));
  INV_X1    g0090(.A(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n216), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G1), .B2(new_n217), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n294), .B1(new_n298), .B2(G50), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT73), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT72), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT71), .B1(new_n301), .B2(new_n201), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT8), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n201), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT71), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n302), .A2(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n217), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n311));
  INV_X1    g0111(.A(G150), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n217), .A2(new_n261), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n296), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n300), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(KEYINPUT9), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n300), .B2(new_n315), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n290), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT10), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n290), .B(new_n322), .C1(new_n317), .C2(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n289), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n288), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n316), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n266), .B2(G20), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n202), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n201), .A2(new_n202), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n206), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  INV_X1    g0141(.A(G159), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n313), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G20), .A2(G33), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT79), .A3(G159), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n331), .B1(new_n338), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n336), .B2(new_n217), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n334), .A2(new_n335), .A3(new_n332), .A4(G20), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(G20), .B1(new_n343), .B2(new_n345), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n348), .A2(new_n296), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n308), .A2(new_n292), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n304), .A2(new_n307), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n298), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n266), .A2(G223), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(G226), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n270), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n285), .A2(G232), .B1(new_n275), .B2(new_n281), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n366), .A2(new_n325), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(G169), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT18), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n360), .A2(new_n373), .A3(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n366), .A2(new_n367), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G200), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(G190), .A3(new_n367), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n355), .A2(new_n359), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n351), .A2(new_n353), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n297), .B1(new_n381), .B2(new_n331), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n383));
  INV_X1    g0183(.A(new_n377), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n259), .B1(new_n366), .B2(new_n367), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT17), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n372), .A2(new_n374), .A3(new_n380), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n330), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n283), .B1(G238), .B2(new_n285), .ZN(new_n391));
  OAI211_X1 g0191(.A(G232), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT76), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n266), .A2(new_n394), .A3(G232), .A4(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n266), .A2(G226), .A3(new_n361), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n393), .A2(new_n395), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT77), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n398), .A2(new_n399), .A3(new_n270), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n398), .B2(new_n270), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n390), .B(new_n391), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n391), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n390), .B1(new_n404), .B2(KEYINPUT78), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(new_n270), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT77), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n398), .A2(new_n399), .A3(new_n270), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT78), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n391), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n403), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G190), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n344), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n230), .B2(new_n309), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n415), .A2(KEYINPUT11), .A3(new_n296), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT12), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n293), .B2(new_n202), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n298), .A2(new_n202), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT11), .B1(new_n415), .B2(new_n296), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n416), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n404), .A2(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n402), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n423), .B1(new_n425), .B2(G200), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n413), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n285), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n282), .B1(new_n428), .B2(new_n231), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT74), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n264), .A2(G232), .B1(new_n336), .B2(G107), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n229), .B2(new_n268), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n270), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n430), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n436), .A2(G179), .ZN(new_n437));
  XOR2_X1   g0237(.A(KEYINPUT8), .B(G58), .Z(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n344), .B1(G20), .B2(G77), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n440), .A2(new_n309), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n297), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n293), .A2(new_n230), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n298), .B2(new_n230), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n436), .A2(new_n327), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n437), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n436), .A2(G200), .ZN(new_n449));
  INV_X1    g0249(.A(G190), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n445), .C1(new_n450), .C2(new_n436), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n389), .A2(new_n427), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n412), .A2(G179), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT14), .B1(new_n425), .B2(G169), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT14), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n457), .B(new_n327), .C1(new_n424), .C2(new_n402), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n423), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n266), .A2(G257), .A3(new_n361), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n266), .A2(G264), .A3(G1698), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n336), .A2(G303), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n270), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n273), .A2(G1), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n281), .A2(G274), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n281), .A2(new_n474), .A3(G270), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n291), .A2(G33), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n292), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n296), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G116), .ZN(new_n481));
  INV_X1    g0281(.A(G116), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n293), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n295), .A2(new_n216), .B1(G20), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n217), .C1(G33), .C2(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT20), .B1(new_n484), .B2(new_n487), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n481), .B(new_n483), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n477), .A2(G169), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT86), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n492), .B(new_n327), .C1(new_n468), .C2(new_n476), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n468), .A2(new_n476), .A3(G179), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n490), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n491), .A2(new_n499), .A3(new_n492), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n490), .B1(new_n477), .B2(G200), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n450), .B2(new_n477), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n494), .A2(new_n498), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n291), .A2(G45), .A3(G274), .ZN(new_n504));
  OAI21_X1  g0304(.A(G250), .B1(new_n273), .B2(G1), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n284), .A2(new_n280), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n507));
  OAI211_X1 g0307(.A(G238), .B(new_n361), .C1(new_n334), .C2(new_n335), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n507), .B(new_n508), .C1(new_n261), .C2(new_n482), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(new_n270), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n327), .ZN(new_n512));
  AOI211_X1 g0312(.A(G179), .B(new_n506), .C1(new_n509), .C2(new_n270), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n217), .B1(new_n396), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G87), .B2(new_n210), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n217), .B(G68), .C1(new_n334), .C2(new_n335), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n309), .B2(new_n486), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n296), .ZN(new_n521));
  INV_X1    g0321(.A(new_n440), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n292), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n480), .A2(new_n522), .ZN(new_n525));
  AND4_X1   g0325(.A1(KEYINPUT85), .A2(new_n521), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n520), .B2(new_n296), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT85), .B1(new_n527), .B2(new_n525), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n512), .B(new_n514), .C1(new_n526), .C2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n479), .A2(new_n530), .A3(new_n296), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n531), .B(new_n523), .C1(new_n520), .C2(new_n296), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n510), .A2(G190), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n533), .C1(new_n259), .C2(new_n510), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n503), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G250), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(new_n361), .C1(new_n334), .C2(new_n335), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n537), .B(new_n485), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT4), .B1(new_n264), .B2(G244), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n270), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n281), .A2(new_n474), .A3(G257), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n471), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n325), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT81), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n313), .B2(new_n230), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n344), .A2(KEYINPUT80), .A3(G77), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT6), .ZN(new_n553));
  AND2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n209), .ZN(new_n555));
  INV_X1    g0355(.A(G107), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n217), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n548), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n551), .ZN(new_n560));
  INV_X1    g0360(.A(new_n557), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n553), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT81), .B(new_n560), .C1(new_n563), .C2(new_n217), .ZN(new_n564));
  OAI21_X1  g0364(.A(G107), .B1(new_n349), .B2(new_n350), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n296), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n293), .A2(new_n486), .ZN(new_n568));
  INV_X1    g0368(.A(new_n480), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(new_n486), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT83), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT83), .B1(new_n542), .B2(new_n544), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n547), .B(new_n572), .C1(new_n575), .C2(G169), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT82), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n567), .B2(new_n571), .ZN(new_n578));
  AOI211_X1 g0378(.A(KEYINPUT82), .B(new_n570), .C1(new_n566), .C2(new_n296), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n545), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT83), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT84), .B1(new_n584), .B2(new_n450), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n545), .A2(G200), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT84), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n575), .A2(new_n587), .A3(G190), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n580), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n536), .A2(new_n576), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n281), .A2(new_n474), .A3(G264), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n281), .A2(new_n474), .A3(KEYINPUT87), .A4(G264), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  OR2_X1    g0396(.A1(G250), .A2(G1698), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(G257), .B2(new_n361), .ZN(new_n598));
  INV_X1    g0398(.A(G294), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n598), .A2(new_n336), .B1(new_n261), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n472), .A2(new_n473), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n504), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n600), .A2(new_n270), .B1(new_n281), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n595), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n596), .B1(new_n595), .B2(new_n603), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n604), .A2(new_n605), .A3(new_n327), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n595), .A2(new_n603), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n325), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT89), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n266), .A2(new_n217), .A3(G87), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT22), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT24), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n261), .A2(new_n482), .A3(G20), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT23), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n217), .B2(G107), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n556), .A2(KEYINPUT23), .A3(G20), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n612), .B1(new_n611), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n296), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n556), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT25), .B1(new_n293), .B2(new_n556), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n569), .A2(new_n556), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n605), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n595), .A2(new_n596), .A3(new_n603), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G169), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT89), .ZN(new_n631));
  INV_X1    g0431(.A(new_n608), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n609), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n450), .B1(new_n604), .B2(new_n605), .ZN(new_n636));
  INV_X1    g0436(.A(new_n607), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(G200), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n611), .A2(new_n617), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT24), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n618), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n625), .B1(new_n641), .B2(new_n296), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n609), .A2(new_n633), .A3(new_n627), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n635), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n463), .A2(new_n590), .A3(new_n646), .ZN(G372));
  NAND2_X1  g0447(.A1(new_n387), .A2(new_n380), .ZN(new_n648));
  INV_X1    g0448(.A(new_n448), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n427), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n460), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n360), .A2(new_n373), .A3(new_n370), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n373), .B1(new_n360), .B2(new_n370), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n324), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n329), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n567), .A2(new_n577), .A3(new_n571), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n510), .B2(new_n259), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n662), .A2(new_n533), .A3(new_n532), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n511), .A2(KEYINPUT91), .A3(G200), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n527), .A2(KEYINPUT85), .A3(new_n525), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n513), .B1(new_n327), .B2(new_n511), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n663), .A2(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n584), .A2(new_n327), .B1(new_n325), .B2(new_n546), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n660), .A2(new_n671), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n576), .B2(new_n535), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n529), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT92), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n674), .A2(new_n675), .A3(new_n678), .A4(new_n529), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n494), .A2(new_n498), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(new_n500), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n627), .B1(new_n606), .B2(new_n608), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n664), .A2(new_n662), .A3(new_n533), .A4(new_n532), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n529), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n638), .B2(new_n642), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n686), .A2(new_n589), .A3(new_n576), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n677), .A2(new_n679), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n657), .B1(new_n463), .B2(new_n688), .ZN(G369));
  NAND3_X1  g0489(.A1(new_n291), .A2(new_n217), .A3(G13), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n490), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n681), .A2(new_n502), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n681), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n695), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n642), .A2(new_n701), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n646), .A2(new_n702), .B1(new_n634), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n682), .A2(new_n695), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n635), .A2(new_n645), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n680), .A2(new_n500), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n701), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n643), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n704), .A2(new_n705), .A3(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n225), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n210), .A2(G87), .A3(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n214), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n635), .A2(new_n681), .A3(new_n645), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n687), .ZN(new_n720));
  INV_X1    g0520(.A(new_n529), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n660), .A2(new_n671), .A3(KEYINPUT26), .A4(new_n673), .ZN(new_n722));
  OAI211_X1 g0522(.A(KEYINPUT95), .B(new_n672), .C1(new_n576), .C2(new_n535), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n672), .B1(new_n576), .B2(new_n535), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n721), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n720), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n701), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  OR3_X1    g0531(.A1(new_n688), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT93), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n510), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n607), .A3(new_n545), .A4(new_n477), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n509), .A2(new_n270), .ZN(new_n738));
  INV_X1    g0538(.A(new_n506), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n600), .A2(new_n270), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n471), .A2(new_n475), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n270), .B2(new_n467), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n741), .A2(new_n743), .A3(G179), .A4(new_n595), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n584), .A2(new_n744), .A3(KEYINPUT30), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n595), .A2(new_n510), .A3(new_n740), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n496), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(new_n575), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n737), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n701), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n735), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n737), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT30), .B1(new_n584), .B2(new_n744), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n575), .A2(new_n746), .A3(new_n748), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n752), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n757), .A2(KEYINPUT93), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT94), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n695), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(KEYINPUT94), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n751), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n536), .A2(new_n576), .A3(new_n589), .A4(new_n701), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n646), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(G330), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n734), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n718), .B1(new_n770), .B2(G1), .ZN(G364));
  NOR2_X1   g0571(.A1(new_n223), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n291), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n713), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n327), .A2(KEYINPUT98), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n217), .B1(KEYINPUT98), .B2(new_n327), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n216), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n217), .A2(new_n325), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n450), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G50), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n217), .A2(G179), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G159), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n785), .A2(new_n786), .B1(new_n791), .B2(KEYINPUT32), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n783), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n794), .A2(new_n202), .B1(new_n795), .B2(new_n530), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n450), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n217), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT99), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G97), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n782), .A2(G190), .A3(new_n259), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n266), .B1(new_n802), .B2(new_n201), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n782), .A2(new_n788), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(G77), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n787), .A2(new_n450), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n791), .A2(KEYINPUT32), .B1(G107), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n797), .A2(new_n801), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n336), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n812), .B(new_n814), .C1(G329), .C2(new_n790), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n784), .A2(G326), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  INV_X1    g0617(.A(new_n795), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n793), .A2(new_n817), .B1(new_n818), .B2(G303), .ZN(new_n819));
  INV_X1    g0619(.A(new_n799), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G294), .B1(new_n808), .B2(G283), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(new_n816), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n781), .B1(new_n810), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n712), .A2(new_n266), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n215), .B2(new_n273), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n254), .B2(new_n273), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n225), .A2(new_n266), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT96), .Z(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G355), .B1(new_n482), .B2(new_n712), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(G13), .A2(G33), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT97), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(G20), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n780), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n776), .B(new_n823), .C1(new_n831), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n834), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n698), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n699), .A2(new_n776), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n698), .A2(G330), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NAND2_X1  g0643(.A1(new_n677), .A2(new_n679), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n683), .A2(new_n687), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n451), .B1(new_n445), .B2(new_n701), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n448), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n649), .A2(new_n701), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n846), .A2(new_n701), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n688), .B2(new_n695), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n775), .B1(new_n854), .B2(new_n768), .ZN(new_n855));
  INV_X1    g0655(.A(new_n768), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n852), .A3(new_n853), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n336), .B1(new_n804), .B2(new_n482), .C1(new_n599), .C2(new_n802), .ZN(new_n859));
  INV_X1    g0659(.A(G283), .ZN(new_n860));
  INV_X1    g0660(.A(G303), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n794), .A2(new_n860), .B1(new_n785), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n859), .B(new_n862), .C1(G107), .C2(new_n818), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n807), .A2(new_n530), .B1(new_n789), .B2(new_n813), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT102), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n863), .A2(new_n801), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n802), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n869), .A2(G143), .B1(new_n805), .B2(G159), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n870), .B1(new_n785), .B2(new_n871), .C1(new_n312), .C2(new_n794), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT34), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n808), .A2(G68), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n336), .B1(new_n790), .B2(G132), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n820), .A2(G58), .B1(new_n818), .B2(G50), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n868), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n781), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  INV_X1    g0683(.A(new_n833), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n780), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT101), .Z(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n776), .B1(new_n887), .B2(new_n230), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n883), .B(new_n888), .C1(new_n851), .C2(new_n833), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT104), .Z(new_n890));
  NOR2_X1   g0690(.A1(new_n858), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  NOR2_X1   g0692(.A1(new_n772), .A2(new_n291), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n733), .A2(new_n462), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n657), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT108), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  INV_X1    g0698(.A(new_n693), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n360), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(KEYINPUT106), .B(new_n693), .C1(new_n355), .C2(new_n359), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n371), .B(new_n378), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n371), .A2(new_n378), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n360), .A2(new_n899), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT106), .B1(new_n383), .B2(new_n693), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n360), .A2(new_n898), .A3(new_n899), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n388), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n908), .A2(KEYINPUT107), .A3(KEYINPUT38), .A4(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT107), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n371), .A2(new_n378), .ZN(new_n914));
  INV_X1    g0714(.A(new_n906), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT37), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n907), .A2(new_n916), .B1(new_n388), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n917), .B2(KEYINPUT38), .ZN(new_n918));
  AND4_X1   g0718(.A1(new_n905), .A2(new_n371), .A3(new_n906), .A4(new_n378), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(KEYINPUT37), .B2(new_n902), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(new_n910), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n387), .A2(new_n380), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n654), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n897), .B(new_n912), .C1(new_n918), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n920), .B2(new_n923), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT39), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n390), .B1(new_n409), .B2(new_n391), .ZN(new_n932));
  OAI21_X1  g0732(.A(G169), .B1(new_n932), .B2(new_n403), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n457), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n425), .A2(KEYINPUT14), .A3(G169), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n935), .B1(G179), .B2(new_n412), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n931), .B1(new_n936), .B2(new_n422), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n459), .A2(KEYINPUT105), .A3(new_n423), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n695), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n852), .A2(new_n849), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n927), .A2(new_n928), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n422), .A2(new_n701), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n413), .B2(new_n426), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n938), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n936), .A2(new_n427), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n942), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n655), .A2(new_n693), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n896), .B(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G330), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n750), .A2(KEYINPUT94), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n757), .A2(new_n761), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT31), .A4(new_n695), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n764), .B(new_n956), .C1(new_n646), .C2(new_n766), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n948), .A2(new_n851), .A3(new_n942), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n918), .A2(new_n925), .ZN(new_n961));
  INV_X1    g0761(.A(new_n912), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n764), .A2(new_n956), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n851), .B1(new_n964), .B2(new_n767), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n963), .A2(new_n966), .A3(KEYINPUT40), .A4(new_n948), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n462), .A2(new_n957), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n953), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n893), .B1(new_n952), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n952), .B2(new_n971), .ZN(new_n973));
  INV_X1    g0773(.A(new_n563), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT35), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT35), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n975), .A2(G116), .A3(new_n218), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT36), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n214), .A2(new_n230), .A3(new_n339), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n786), .B2(G68), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n223), .A2(G1), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n973), .B(new_n978), .C1(new_n980), .C2(new_n981), .ZN(G367));
  OAI211_X1 g0782(.A(new_n589), .B(new_n576), .C1(new_n580), .C2(new_n701), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n660), .A2(new_n673), .A3(new_n695), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n710), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n576), .B1(new_n985), .B2(new_n706), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n701), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n671), .B1(new_n532), .B2(new_n701), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n529), .A2(new_n532), .A3(new_n701), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n990), .A2(new_n991), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT43), .B1(new_n995), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n704), .A2(new_n985), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n999), .A2(new_n1000), .B1(new_n704), .B2(new_n985), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n713), .B(KEYINPUT41), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n710), .A2(new_n705), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n985), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT44), .Z(new_n1008));
  NOR2_X1   g0808(.A1(new_n1006), .A2(new_n985), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1011), .A2(new_n700), .A3(new_n703), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n710), .B1(new_n703), .B2(new_n709), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n699), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n769), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1008), .A2(new_n704), .A3(new_n1010), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1005), .B1(new_n1017), .B2(new_n770), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1003), .B(new_n1004), .C1(new_n774), .C2(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n249), .A2(new_n824), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n835), .B1(new_n225), .B2(new_n440), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n775), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n266), .B1(new_n802), .B2(new_n312), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n807), .A2(new_n230), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G143), .B2(new_n784), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n342), .B2(new_n794), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(G50), .C2(new_n805), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n818), .A2(G58), .B1(new_n790), .B2(G137), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT111), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n800), .A2(G68), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(KEYINPUT111), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n793), .A2(G294), .B1(new_n808), .B2(G97), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n556), .B2(new_n799), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n785), .A2(new_n813), .B1(new_n861), .B2(new_n802), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(KEYINPUT110), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n336), .B1(new_n789), .B2(new_n1037), .C1(new_n860), .C2(new_n804), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n818), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT46), .B1(new_n818), .B2(G116), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1036), .B(new_n1041), .C1(KEYINPUT110), .C2(new_n1035), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1032), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1022), .B1(new_n1044), .B2(new_n780), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n837), .B2(new_n996), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1019), .A2(new_n1046), .ZN(G387));
  NOR2_X1   g0847(.A1(new_n1015), .A2(new_n714), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1014), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n770), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n703), .A2(new_n837), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n715), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n829), .A2(new_n1052), .B1(new_n556), .B2(new_n712), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n245), .A2(new_n273), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n438), .A2(new_n786), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n715), .B(new_n273), .C1(new_n202), .C2(new_n230), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n824), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1059), .A2(new_n835), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n785), .A2(new_n342), .B1(new_n807), .B2(new_n486), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n869), .A2(G50), .B1(new_n790), .B2(G150), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n266), .C1(new_n202), .C2(new_n804), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(G77), .C2(new_n818), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n800), .A2(new_n522), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n308), .C2(new_n794), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT112), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n869), .A2(G317), .B1(new_n805), .B2(G303), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT113), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n793), .A2(G311), .B1(new_n784), .B2(G322), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n799), .A2(new_n860), .B1(new_n795), .B2(new_n599), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT49), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(KEYINPUT49), .A3(new_n1076), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n266), .B1(new_n790), .B2(G326), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n482), .C2(new_n807), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1067), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n776), .B(new_n1060), .C1(new_n1081), .C2(new_n780), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1049), .A2(new_n774), .B1(new_n1051), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1050), .A2(new_n1083), .ZN(G393));
  NAND2_X1  g0884(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(new_n773), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n985), .A2(new_n834), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n835), .B1(new_n486), .B2(new_n225), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n825), .A2(new_n257), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n775), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n785), .A2(new_n312), .B1(new_n342), .B2(new_n802), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT114), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n336), .B1(new_n790), .B2(G143), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n202), .B2(new_n795), .C1(new_n530), .C2(new_n807), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1092), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1093), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n793), .A2(G50), .B1(new_n805), .B2(new_n438), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n800), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1097), .B(new_n1098), .C1(new_n230), .C2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G317), .A2(new_n784), .B1(new_n869), .B2(G311), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n794), .A2(new_n861), .B1(new_n807), .B2(new_n556), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n336), .B1(new_n789), .B2(new_n811), .C1(new_n599), .C2(new_n804), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n799), .A2(new_n482), .B1(new_n795), .B2(new_n860), .ZN(new_n1105));
  OR3_X1    g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1096), .A2(new_n1100), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1090), .B1(new_n1107), .B2(new_n780), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1086), .B1(new_n1087), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1085), .B1(new_n769), .B2(new_n1014), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(new_n713), .A3(new_n1017), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(G390));
  AOI21_X1  g0912(.A(new_n948), .B1(new_n966), .B2(G330), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n848), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n849), .B1(new_n730), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n851), .C1(new_n765), .C2(new_n767), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT115), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n1119), .A3(new_n948), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n945), .A2(new_n947), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT115), .B1(new_n1121), .B2(new_n1117), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n966), .A2(G330), .A3(new_n948), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n948), .B2(new_n1118), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n941), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n462), .A2(G330), .A3(new_n957), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n894), .A2(new_n657), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1125), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n688), .A2(new_n695), .A3(new_n850), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n849), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n948), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n939), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n930), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n927), .B(new_n913), .C1(KEYINPUT38), .C2(new_n917), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1139), .A3(new_n912), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1115), .B2(new_n948), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1133), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n926), .A2(new_n929), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n852), .A2(new_n849), .B1(new_n945), .B2(new_n947), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n939), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n695), .B1(new_n720), .B2(new_n728), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1135), .B1(new_n1146), .B2(new_n848), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1137), .B(new_n963), .C1(new_n1147), .C2(new_n1121), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1123), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n714), .B1(new_n1132), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1132), .B2(new_n1150), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1143), .A2(new_n884), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n775), .B1(new_n886), .B2(new_n357), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n795), .A2(new_n312), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1099), .B2(new_n342), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n784), .A2(G128), .B1(new_n808), .B2(G50), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n871), .B2(new_n794), .ZN(new_n1159));
  INV_X1    g0959(.A(G132), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n266), .B1(new_n802), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n804), .A2(new_n1162), .B1(new_n789), .B2(new_n1163), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1157), .A2(new_n1159), .A3(new_n1161), .A4(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT116), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(KEYINPUT116), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n784), .A2(G283), .B1(new_n805), .B2(G97), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n556), .B2(new_n794), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n336), .B1(new_n795), .B2(new_n530), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT118), .Z(new_n1172));
  OAI221_X1 g0972(.A(new_n876), .B1(new_n482), .B2(new_n802), .C1(new_n599), .C2(new_n789), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G77), .B2(new_n800), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1166), .A2(new_n1167), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1154), .B1(new_n1176), .B2(new_n780), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1153), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1150), .B2(new_n773), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1152), .B1(new_n1180), .B2(new_n1181), .ZN(G378));
  AOI21_X1  g0982(.A(new_n693), .B1(new_n300), .B2(new_n315), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n330), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT123), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1183), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n324), .A2(new_n329), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n324), .B2(new_n329), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n329), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1190), .B(new_n1183), .C1(new_n321), .C2(new_n323), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT123), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1193));
  AND3_X1   g0993(.A1(new_n1188), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND4_X1   g0996(.A1(G330), .A2(new_n960), .A3(new_n967), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n965), .B1(new_n945), .B2(new_n947), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n961), .A2(new_n959), .A3(new_n962), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n953), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1196), .B1(new_n1200), .B2(new_n960), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n951), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT124), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n960), .A2(G330), .A3(new_n967), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1196), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n940), .A2(new_n949), .A3(new_n950), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1200), .A2(new_n960), .A3(new_n1196), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1203), .A3(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1123), .A2(new_n1116), .B1(new_n1126), .B2(new_n941), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1131), .B1(new_n1150), .B2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1206), .A2(new_n1207), .A3(KEYINPUT124), .A4(new_n1208), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1202), .B2(new_n1209), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n714), .B1(new_n1217), .B2(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1210), .A2(new_n774), .A3(new_n1213), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n885), .A2(new_n786), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(new_n775), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G41), .B(new_n266), .C1(new_n790), .C2(G283), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n201), .B2(new_n807), .C1(new_n230), .C2(new_n795), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT121), .Z(new_n1225));
  AOI22_X1  g1025(.A1(new_n869), .A2(G107), .B1(new_n805), .B2(new_n522), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n785), .B2(new_n482), .C1(new_n486), .C2(new_n794), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G68), .B2(new_n800), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(KEYINPUT58), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(G33), .A2(G41), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT120), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n786), .C1(G41), .C2(new_n266), .ZN(new_n1235));
  INV_X1    g1035(.A(G128), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n802), .A2(new_n1236), .B1(new_n804), .B2(new_n871), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G132), .B2(new_n793), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1162), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n784), .A2(G125), .B1(new_n818), .B2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(new_n1099), .C2(new_n312), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n807), .A2(new_n342), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(KEYINPUT122), .B(G124), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1234), .B(new_n1244), .C1(new_n790), .C2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1242), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  AND4_X1   g1047(.A1(new_n1229), .A2(new_n1232), .A3(new_n1235), .A4(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1222), .B1(new_n781), .B2(new_n1248), .C1(new_n1196), .C2(new_n833), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1220), .A2(KEYINPUT125), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT125), .B1(new_n1220), .B2(new_n1249), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1219), .B1(new_n1250), .B2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1211), .A2(new_n1130), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1005), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1132), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n802), .A2(new_n860), .B1(new_n804), .B2(new_n556), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n266), .B(new_n1256), .C1(G303), .C2(new_n790), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1024), .B1(G116), .B2(new_n793), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n784), .A2(G294), .B1(new_n818), .B2(G97), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1257), .A2(new_n1065), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n804), .A2(new_n312), .B1(new_n789), .B2(new_n1236), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n336), .B(new_n1261), .C1(G137), .C2(new_n869), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n800), .A2(G50), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n784), .A2(G132), .B1(new_n808), .B2(G58), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n793), .A2(new_n1239), .B1(new_n818), .B2(G159), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n781), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n776), .B(new_n1267), .C1(new_n202), .C2(new_n887), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n948), .B2(new_n833), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1211), .B2(new_n773), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1255), .A2(new_n1271), .ZN(G381));
  NAND3_X1  g1072(.A1(new_n1050), .A2(new_n842), .A3(new_n1083), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1179), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1152), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  OR4_X1    g1077(.A1(G387), .A2(new_n1274), .A3(G375), .A4(new_n1277), .ZN(G407));
  NAND2_X1  g1078(.A1(new_n694), .A2(G213), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G407), .B(G213), .C1(G375), .C2(new_n1281), .ZN(G409));
  NAND2_X1  g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1273), .ZN(new_n1285));
  OR3_X1    g1085(.A1(new_n1284), .A2(KEYINPUT126), .A3(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1019), .B2(new_n1046), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1019), .A2(G390), .A3(new_n1046), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1291), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1293), .B2(new_n1289), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1219), .B(G378), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1202), .A2(new_n1209), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n1249), .B1(new_n773), .B2(new_n1298), .C1(new_n1214), .C2(new_n1005), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1276), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1253), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1211), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n713), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(G384), .A3(new_n1271), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n713), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1303), .B2(new_n1253), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n891), .B1(new_n1309), .B2(new_n1270), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1301), .A2(new_n1302), .A3(new_n1279), .A4(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1280), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1280), .A2(G2897), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1307), .A2(new_n1310), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1313), .B(new_n1314), .C1(new_n1315), .C2(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1315), .B2(new_n1312), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1296), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1315), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1325), .B2(new_n1311), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1312), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1328), .A3(new_n1295), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1323), .A2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1276), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1311), .A3(new_n1297), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1311), .B1(new_n1332), .B2(new_n1297), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1295), .ZN(G402));
endmodule


