

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794;

  XNOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n361) );
  XOR2_X1 U383 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n362) );
  XNOR2_X1 U384 ( .A(KEYINPUT59), .B(n675), .ZN(n363) );
  AND2_X1 U385 ( .A1(n442), .A2(n385), .ZN(n364) );
  NOR2_X2 U386 ( .A1(n733), .A2(n619), .ZN(n622) );
  OR2_X2 U387 ( .A1(n717), .A2(n635), .ZN(n631) );
  XNOR2_X2 U388 ( .A(n481), .B(n480), .ZN(n569) );
  NOR2_X2 U389 ( .A1(n676), .A2(n794), .ZN(n634) );
  XNOR2_X2 U390 ( .A(n632), .B(n633), .ZN(n676) );
  AND2_X1 U391 ( .A1(n370), .A2(n368), .ZN(n367) );
  AND2_X1 U392 ( .A1(n369), .A2(n605), .ZN(n368) );
  INV_X1 U393 ( .A(n572), .ZN(n549) );
  INV_X1 U394 ( .A(G475), .ZN(n416) );
  NOR2_X1 U395 ( .A1(n755), .A2(n754), .ZN(n757) );
  XNOR2_X1 U396 ( .A(n378), .B(n363), .ZN(n377) );
  NAND2_X1 U397 ( .A1(n409), .A2(n410), .ZN(n378) );
  NAND2_X1 U398 ( .A1(n373), .A2(n375), .ZN(n374) );
  NAND2_X1 U399 ( .A1(n438), .A2(n440), .ZN(n375) );
  AND2_X1 U400 ( .A1(n364), .A2(n443), .ZN(n373) );
  NAND2_X1 U401 ( .A1(n367), .A2(n366), .ZN(n544) );
  NAND2_X1 U402 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U403 ( .A(n403), .B(n387), .ZN(n713) );
  NOR2_X1 U404 ( .A1(n380), .A2(n513), .ZN(n371) );
  NAND2_X1 U405 ( .A1(n425), .A2(n422), .ZN(n750) );
  BUF_X1 U406 ( .A(n592), .Z(n391) );
  XNOR2_X1 U407 ( .A(n478), .B(n477), .ZN(n589) );
  XNOR2_X1 U408 ( .A(n517), .B(n463), .ZN(n662) );
  INV_X1 U409 ( .A(n701), .ZN(n365) );
  INV_X1 U410 ( .A(n776), .ZN(n455) );
  XNOR2_X1 U411 ( .A(n498), .B(n462), .ZN(n517) );
  XOR2_X1 U412 ( .A(KEYINPUT75), .B(KEYINPUT34), .Z(n513) );
  NAND2_X1 U413 ( .A1(n713), .A2(n513), .ZN(n366) );
  NAND2_X1 U414 ( .A1(n380), .A2(n513), .ZN(n369) );
  INV_X1 U415 ( .A(n713), .ZN(n372) );
  XNOR2_X2 U416 ( .A(n374), .B(n361), .ZN(n649) );
  XNOR2_X1 U417 ( .A(n376), .B(n362), .ZN(G60) );
  NAND2_X1 U418 ( .A1(n377), .A2(n365), .ZN(n376) );
  INV_X1 U419 ( .A(n439), .ZN(n379) );
  INV_X1 U420 ( .A(n549), .ZN(n380) );
  XNOR2_X1 U421 ( .A(n556), .B(n555), .ZN(n678) );
  XNOR2_X1 U422 ( .A(n512), .B(KEYINPUT0), .ZN(n572) );
  NOR2_X1 U423 ( .A1(n649), .A2(n661), .ZN(n381) );
  XNOR2_X1 U424 ( .A(n610), .B(n461), .ZN(n382) );
  NOR2_X1 U425 ( .A1(n649), .A2(n661), .ZN(n703) );
  XNOR2_X1 U426 ( .A(n610), .B(n461), .ZN(n552) );
  XNOR2_X1 U427 ( .A(n399), .B(n483), .ZN(n496) );
  XNOR2_X1 U428 ( .A(G119), .B(G116), .ZN(n483) );
  XNOR2_X1 U429 ( .A(n484), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U430 ( .A(G113), .B(KEYINPUT71), .ZN(n484) );
  NOR2_X1 U431 ( .A1(n715), .A2(n600), .ZN(n601) );
  AND2_X1 U432 ( .A1(n617), .A2(n616), .ZN(n421) );
  XOR2_X1 U433 ( .A(G137), .B(KEYINPUT5), .Z(n487) );
  XNOR2_X1 U434 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n462) );
  XNOR2_X1 U435 ( .A(G134), .B(G131), .ZN(n663) );
  INV_X1 U436 ( .A(KEYINPUT1), .ZN(n461) );
  XNOR2_X1 U437 ( .A(n407), .B(n465), .ZN(n406) );
  XNOR2_X1 U438 ( .A(n467), .B(n466), .ZN(n407) );
  XNOR2_X1 U439 ( .A(G128), .B(G119), .ZN(n464) );
  NAND2_X1 U440 ( .A1(n383), .A2(n646), .ZN(n436) );
  XNOR2_X1 U441 ( .A(n501), .B(n498), .ZN(n419) );
  XNOR2_X1 U442 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n500) );
  XNOR2_X1 U443 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n499) );
  XNOR2_X1 U444 ( .A(n496), .B(n495), .ZN(n778) );
  XNOR2_X1 U445 ( .A(KEYINPUT16), .B(G122), .ZN(n494) );
  XNOR2_X1 U446 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n550) );
  NOR2_X1 U447 ( .A1(n720), .A2(n547), .ZN(n548) );
  XNOR2_X1 U448 ( .A(n773), .B(KEYINPUT91), .ZN(n617) );
  XNOR2_X1 U449 ( .A(G110), .B(KEYINPUT23), .ZN(n466) );
  XOR2_X1 U450 ( .A(G131), .B(KEYINPUT103), .Z(n516) );
  XNOR2_X1 U451 ( .A(G143), .B(G113), .ZN(n519) );
  XOR2_X1 U452 ( .A(G122), .B(G104), .Z(n520) );
  NAND2_X1 U453 ( .A1(n383), .A2(n388), .ZN(n437) );
  NOR2_X1 U454 ( .A1(n720), .A2(KEYINPUT41), .ZN(n423) );
  NAND2_X1 U455 ( .A1(n622), .A2(n719), .ZN(n623) );
  INV_X1 U456 ( .A(G902), .ZN(n583) );
  XNOR2_X1 U457 ( .A(n400), .B(n496), .ZN(n490) );
  XNOR2_X1 U458 ( .A(n488), .B(n485), .ZN(n400) );
  INV_X1 U459 ( .A(G953), .ZN(n783) );
  INV_X1 U460 ( .A(G128), .ZN(n451) );
  XNOR2_X1 U461 ( .A(G116), .B(G134), .ZN(n530) );
  AND2_X1 U462 ( .A1(n427), .A2(n426), .ZN(n425) );
  NAND2_X1 U463 ( .A1(n424), .A2(n423), .ZN(n422) );
  NAND2_X1 U464 ( .A1(n720), .A2(KEYINPUT41), .ZN(n426) );
  NAND2_X1 U465 ( .A1(n402), .A2(n401), .ZN(n636) );
  XNOR2_X1 U466 ( .A(n391), .B(n386), .ZN(n392) );
  INV_X1 U467 ( .A(G469), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n592), .B(n386), .ZN(n511) );
  INV_X1 U469 ( .A(G472), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n470), .B(n405), .ZN(n694) );
  XNOR2_X1 U471 ( .A(n778), .B(n418), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n419), .B(n497), .ZN(n418) );
  INV_X1 U473 ( .A(G210), .ZN(n412) );
  NOR2_X1 U474 ( .A1(n668), .A2(G952), .ZN(n701) );
  INV_X1 U475 ( .A(G140), .ZN(n657) );
  XNOR2_X1 U476 ( .A(n629), .B(n628), .ZN(n794) );
  AND2_X1 U477 ( .A1(n397), .A2(n594), .ZN(n773) );
  XNOR2_X1 U478 ( .A(n398), .B(KEYINPUT36), .ZN(n397) );
  NOR2_X1 U479 ( .A1(n593), .A2(n391), .ZN(n398) );
  XNOR2_X1 U480 ( .A(n636), .B(KEYINPUT114), .ZN(n593) );
  NAND2_X1 U481 ( .A1(n648), .A2(KEYINPUT67), .ZN(n383) );
  XNOR2_X1 U482 ( .A(n553), .B(n493), .ZN(n591) );
  INV_X1 U483 ( .A(n591), .ZN(n401) );
  AND2_X1 U484 ( .A1(n599), .A2(n610), .ZN(n384) );
  AND2_X1 U485 ( .A1(n582), .A2(n659), .ZN(n385) );
  XOR2_X1 U486 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n386) );
  XNOR2_X1 U487 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n387) );
  OR2_X1 U488 ( .A1(n645), .A2(KEYINPUT67), .ZN(n388) );
  XOR2_X1 U489 ( .A(KEYINPUT90), .B(KEYINPUT48), .Z(n389) );
  XNOR2_X1 U490 ( .A(G902), .B(KEYINPUT15), .ZN(n646) );
  XNOR2_X1 U491 ( .A(n390), .B(n694), .ZN(n695) );
  AND2_X1 U492 ( .A1(n696), .A2(G217), .ZN(n390) );
  NOR2_X1 U493 ( .A1(n434), .A2(n710), .ZN(n696) );
  NOR2_X1 U494 ( .A1(n441), .A2(n439), .ZN(n438) );
  BUF_X1 U495 ( .A(n589), .Z(n558) );
  OR2_X2 U496 ( .A1(n621), .A2(n635), .ZN(n592) );
  AND2_X1 U497 ( .A1(n615), .A2(n450), .ZN(n616) );
  NOR2_X1 U498 ( .A1(n627), .A2(n595), .ZN(n402) );
  XNOR2_X1 U499 ( .A(n662), .B(n406), .ZN(n405) );
  XNOR2_X2 U500 ( .A(n394), .B(n393), .ZN(n610) );
  NOR2_X1 U501 ( .A1(n698), .A2(G902), .ZN(n394) );
  NOR2_X1 U502 ( .A1(n710), .A2(n412), .ZN(n411) );
  NOR2_X1 U503 ( .A1(n710), .A2(n414), .ZN(n413) );
  NAND2_X1 U504 ( .A1(n415), .A2(n411), .ZN(n683) );
  NAND2_X1 U505 ( .A1(n415), .A2(n413), .ZN(n689) );
  OR2_X2 U506 ( .A1(n703), .A2(n437), .ZN(n435) );
  NOR2_X1 U507 ( .A1(n684), .A2(n701), .ZN(n685) );
  NOR2_X1 U508 ( .A1(n690), .A2(n701), .ZN(n692) );
  NAND2_X1 U509 ( .A1(n421), .A2(n420), .ZN(n396) );
  XNOR2_X2 U510 ( .A(n650), .B(n644), .ZN(n661) );
  NAND2_X1 U511 ( .A1(n395), .A2(n643), .ZN(n650) );
  XNOR2_X1 U512 ( .A(n396), .B(n389), .ZN(n395) );
  XNOR2_X2 U513 ( .A(n492), .B(n491), .ZN(n553) );
  NAND2_X1 U514 ( .A1(n404), .A2(n401), .ZN(n403) );
  XNOR2_X1 U515 ( .A(n566), .B(KEYINPUT110), .ZN(n404) );
  OR2_X2 U516 ( .A1(n431), .A2(n428), .ZN(n566) );
  XNOR2_X1 U517 ( .A(n408), .B(n417), .ZN(n681) );
  XNOR2_X1 U518 ( .A(n408), .B(n460), .ZN(n698) );
  XNOR2_X2 U519 ( .A(n489), .B(n455), .ZN(n408) );
  NOR2_X1 U520 ( .A1(n710), .A2(n416), .ZN(n409) );
  INV_X1 U521 ( .A(n434), .ZN(n410) );
  INV_X1 U522 ( .A(n434), .ZN(n415) );
  NAND2_X1 U523 ( .A1(n384), .A2(n392), .ZN(n763) );
  NOR2_X2 U524 ( .A1(n782), .A2(n652), .ZN(n710) );
  XNOR2_X2 U525 ( .A(n667), .B(n453), .ZN(n489) );
  XNOR2_X2 U526 ( .A(n535), .B(KEYINPUT4), .ZN(n667) );
  XNOR2_X1 U527 ( .A(n634), .B(KEYINPUT46), .ZN(n420) );
  NAND2_X1 U528 ( .A1(n750), .A2(n384), .ZN(n632) );
  INV_X1 U529 ( .A(n716), .ZN(n424) );
  NAND2_X1 U530 ( .A1(n716), .A2(KEYINPUT41), .ZN(n427) );
  XNOR2_X2 U531 ( .A(n631), .B(n630), .ZN(n716) );
  NAND2_X1 U532 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U533 ( .A1(n569), .A2(n482), .ZN(n429) );
  NAND2_X1 U534 ( .A1(n552), .A2(n482), .ZN(n430) );
  NOR2_X1 U535 ( .A1(n382), .A2(n432), .ZN(n431) );
  NAND2_X1 U536 ( .A1(n433), .A2(KEYINPUT78), .ZN(n432) );
  INV_X1 U537 ( .A(n569), .ZN(n433) );
  NAND2_X2 U538 ( .A1(n435), .A2(n436), .ZN(n434) );
  INV_X1 U539 ( .A(n678), .ZN(n439) );
  INV_X1 U540 ( .A(n693), .ZN(n440) );
  XNOR2_X2 U541 ( .A(n544), .B(KEYINPUT35), .ZN(n693) );
  NAND2_X1 U542 ( .A1(n678), .A2(n660), .ZN(n445) );
  NAND2_X1 U543 ( .A1(n660), .A2(n565), .ZN(n441) );
  NAND2_X1 U544 ( .A1(n445), .A2(n444), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n693), .A2(n444), .ZN(n443) );
  INV_X1 U546 ( .A(n565), .ZN(n444) );
  AND2_X1 U547 ( .A1(n655), .A2(n365), .ZN(G63) );
  AND2_X1 U548 ( .A1(n479), .A2(G221), .ZN(n447) );
  AND2_X1 U549 ( .A1(n746), .A2(n510), .ZN(n448) );
  NAND2_X1 U550 ( .A1(n656), .A2(n613), .ZN(n449) );
  NOR2_X1 U551 ( .A1(n614), .A2(n449), .ZN(n450) );
  NAND2_X1 U552 ( .A1(n511), .A2(n448), .ZN(n512) );
  NOR2_X1 U553 ( .A1(n624), .A2(n623), .ZN(n626) );
  INV_X1 U554 ( .A(KEYINPUT40), .ZN(n628) );
  INV_X1 U555 ( .A(KEYINPUT109), .ZN(n555) );
  XNOR2_X2 U556 ( .A(G143), .B(KEYINPUT84), .ZN(n452) );
  XNOR2_X2 U557 ( .A(n452), .B(n451), .ZN(n535) );
  XNOR2_X1 U558 ( .A(KEYINPUT68), .B(G101), .ZN(n453) );
  XNOR2_X1 U559 ( .A(G110), .B(G107), .ZN(n454) );
  XNOR2_X1 U560 ( .A(n454), .B(G104), .ZN(n776) );
  XNOR2_X1 U561 ( .A(n663), .B(G146), .ZN(n485) );
  XNOR2_X1 U562 ( .A(n657), .B(G137), .ZN(n463) );
  XNOR2_X1 U563 ( .A(n463), .B(KEYINPUT82), .ZN(n458) );
  INV_X1 U564 ( .A(KEYINPUT64), .ZN(n456) );
  XNOR2_X2 U565 ( .A(n456), .B(G953), .ZN(n668) );
  NAND2_X1 U566 ( .A1(n668), .A2(G227), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U568 ( .A(n485), .B(n459), .ZN(n460) );
  XNOR2_X2 U569 ( .A(G125), .B(G146), .ZN(n498) );
  XNOR2_X1 U570 ( .A(KEYINPUT97), .B(n464), .ZN(n465) );
  XOR2_X1 U571 ( .A(KEYINPUT24), .B(KEYINPUT72), .Z(n467) );
  NAND2_X1 U572 ( .A1(n668), .A2(G234), .ZN(n468) );
  XNOR2_X1 U573 ( .A(n468), .B(KEYINPUT8), .ZN(n538) );
  INV_X1 U574 ( .A(G221), .ZN(n469) );
  OR2_X1 U575 ( .A1(n538), .A2(n469), .ZN(n470) );
  NAND2_X1 U576 ( .A1(n694), .A2(n583), .ZN(n478) );
  NAND2_X1 U577 ( .A1(n646), .A2(G234), .ZN(n471) );
  XNOR2_X1 U578 ( .A(n471), .B(KEYINPUT20), .ZN(n472) );
  XNOR2_X1 U579 ( .A(KEYINPUT98), .B(n472), .ZN(n479) );
  AND2_X1 U580 ( .A1(n479), .A2(G217), .ZN(n476) );
  XNOR2_X1 U581 ( .A(KEYINPUT81), .B(KEYINPUT99), .ZN(n474) );
  XNOR2_X1 U582 ( .A(KEYINPUT25), .B(KEYINPUT80), .ZN(n473) );
  XNOR2_X1 U583 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U584 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U585 ( .A(KEYINPUT21), .B(n447), .ZN(n727) );
  XNOR2_X1 U586 ( .A(n727), .B(KEYINPUT100), .ZN(n546) );
  NAND2_X1 U587 ( .A1(n589), .A2(n546), .ZN(n481) );
  INV_X1 U588 ( .A(KEYINPUT69), .ZN(n480) );
  INV_X1 U589 ( .A(KEYINPUT78), .ZN(n482) );
  NOR2_X1 U590 ( .A1(G953), .A2(G237), .ZN(n514) );
  NAND2_X1 U591 ( .A1(n514), .A2(G210), .ZN(n486) );
  XNOR2_X1 U592 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U593 ( .A(n489), .B(n490), .ZN(n687) );
  NAND2_X1 U594 ( .A1(n687), .A2(n583), .ZN(n492) );
  XOR2_X1 U595 ( .A(G472), .B(KEYINPUT101), .Z(n491) );
  XOR2_X1 U596 ( .A(KEYINPUT107), .B(KEYINPUT6), .Z(n493) );
  XNOR2_X1 U597 ( .A(n494), .B(KEYINPUT76), .ZN(n495) );
  NAND2_X1 U598 ( .A1(n668), .A2(G224), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U600 ( .A(n646), .ZN(n647) );
  NOR2_X1 U601 ( .A1(n681), .A2(n647), .ZN(n505) );
  INV_X1 U602 ( .A(G237), .ZN(n502) );
  NAND2_X1 U603 ( .A1(n583), .A2(n502), .ZN(n506) );
  NAND2_X1 U604 ( .A1(n506), .A2(G210), .ZN(n503) );
  XOR2_X1 U605 ( .A(n503), .B(KEYINPUT96), .Z(n504) );
  XNOR2_X2 U606 ( .A(n505), .B(n504), .ZN(n621) );
  NAND2_X1 U607 ( .A1(n506), .A2(G214), .ZN(n718) );
  INV_X1 U608 ( .A(n718), .ZN(n635) );
  NAND2_X1 U609 ( .A1(G237), .A2(G234), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n507), .B(KEYINPUT14), .ZN(n746) );
  INV_X1 U611 ( .A(G898), .ZN(n779) );
  AND2_X1 U612 ( .A1(n779), .A2(G902), .ZN(n508) );
  NAND2_X1 U613 ( .A1(n508), .A2(G953), .ZN(n509) );
  NAND2_X1 U614 ( .A1(n783), .A2(G952), .ZN(n587) );
  NAND2_X1 U615 ( .A1(n509), .A2(n587), .ZN(n510) );
  NAND2_X1 U616 ( .A1(G214), .A2(n514), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U618 ( .A(n518), .B(n517), .Z(n526) );
  XNOR2_X1 U619 ( .A(n520), .B(n519), .ZN(n524) );
  XOR2_X1 U620 ( .A(KEYINPUT104), .B(KEYINPUT11), .Z(n522) );
  XNOR2_X1 U621 ( .A(G140), .B(KEYINPUT12), .ZN(n521) );
  XNOR2_X1 U622 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U623 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U624 ( .A(n526), .B(n525), .ZN(n675) );
  NOR2_X1 U625 ( .A1(G902), .A2(n675), .ZN(n528) );
  XNOR2_X1 U626 ( .A(KEYINPUT105), .B(KEYINPUT13), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n529), .B(G475), .ZN(n574) );
  INV_X1 U629 ( .A(n574), .ZN(n542) );
  XNOR2_X1 U630 ( .A(n530), .B(G107), .ZN(n534) );
  XOR2_X1 U631 ( .A(KEYINPUT9), .B(KEYINPUT106), .Z(n532) );
  XNOR2_X1 U632 ( .A(G122), .B(KEYINPUT7), .ZN(n531) );
  XNOR2_X1 U633 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U634 ( .A(n534), .B(n533), .Z(n536) );
  XNOR2_X1 U635 ( .A(n535), .B(n536), .ZN(n540) );
  INV_X1 U636 ( .A(G217), .ZN(n537) );
  OR2_X1 U637 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n540), .B(n539), .ZN(n653) );
  NAND2_X1 U639 ( .A1(n653), .A2(n583), .ZN(n541) );
  XNOR2_X1 U640 ( .A(n541), .B(G478), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n542), .A2(n573), .ZN(n543) );
  XNOR2_X1 U642 ( .A(n543), .B(KEYINPUT111), .ZN(n605) );
  INV_X1 U643 ( .A(n573), .ZN(n545) );
  NAND2_X1 U644 ( .A1(n574), .A2(n545), .ZN(n720) );
  INV_X1 U645 ( .A(n546), .ZN(n547) );
  NAND2_X1 U646 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U647 ( .A(n551), .B(n550), .ZN(n557) );
  INV_X1 U648 ( .A(n382), .ZN(n594) );
  NOR2_X1 U649 ( .A1(n557), .A2(n594), .ZN(n581) );
  NOR2_X1 U650 ( .A1(n553), .A2(n558), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n581), .A2(n554), .ZN(n556) );
  INV_X1 U652 ( .A(n557), .ZN(n562) );
  XOR2_X1 U653 ( .A(KEYINPUT108), .B(n558), .Z(n729) );
  NAND2_X1 U654 ( .A1(n594), .A2(n729), .ZN(n560) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT83), .ZN(n559) );
  NOR2_X1 U656 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U657 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U658 ( .A(n563), .B(KEYINPUT32), .ZN(n660) );
  INV_X1 U659 ( .A(KEYINPUT74), .ZN(n564) );
  NOR2_X1 U660 ( .A1(n564), .A2(KEYINPUT44), .ZN(n565) );
  NAND2_X1 U661 ( .A1(n566), .A2(n553), .ZN(n737) );
  NOR2_X1 U662 ( .A1(n572), .A2(n737), .ZN(n568) );
  XOR2_X1 U663 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n567) );
  XNOR2_X1 U664 ( .A(n568), .B(n567), .ZN(n771) );
  BUF_X2 U665 ( .A(n569), .Z(n733) );
  NOR2_X1 U666 ( .A1(n733), .A2(n553), .ZN(n570) );
  NAND2_X1 U667 ( .A1(n570), .A2(n610), .ZN(n571) );
  NOR2_X1 U668 ( .A1(n380), .A2(n571), .ZN(n759) );
  NOR2_X1 U669 ( .A1(n771), .A2(n759), .ZN(n576) );
  AND2_X1 U670 ( .A1(n574), .A2(n573), .ZN(n770) );
  INV_X1 U671 ( .A(n770), .ZN(n575) );
  OR2_X1 U672 ( .A1(n574), .A2(n573), .ZN(n627) );
  AND2_X1 U673 ( .A1(n575), .A2(n627), .ZN(n715) );
  NOR2_X1 U674 ( .A1(n576), .A2(n715), .ZN(n579) );
  INV_X1 U675 ( .A(KEYINPUT44), .ZN(n577) );
  NOR2_X1 U676 ( .A1(n577), .A2(KEYINPUT74), .ZN(n578) );
  NOR2_X1 U677 ( .A1(n579), .A2(n578), .ZN(n582) );
  NOR2_X1 U678 ( .A1(n401), .A2(n729), .ZN(n580) );
  NAND2_X1 U679 ( .A1(n581), .A2(n580), .ZN(n659) );
  NOR2_X1 U680 ( .A1(G900), .A2(n583), .ZN(n585) );
  INV_X1 U681 ( .A(n668), .ZN(n584) );
  NAND2_X1 U682 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U683 ( .A1(n587), .A2(n586), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n727), .A2(n603), .ZN(n588) );
  NOR2_X1 U685 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U686 ( .A1(n746), .A2(n590), .ZN(n595) );
  INV_X1 U687 ( .A(n595), .ZN(n596) );
  NAND2_X1 U688 ( .A1(n553), .A2(n596), .ZN(n598) );
  INV_X1 U689 ( .A(KEYINPUT28), .ZN(n597) );
  XNOR2_X1 U690 ( .A(n598), .B(n597), .ZN(n599) );
  OR2_X1 U691 ( .A1(n763), .A2(KEYINPUT47), .ZN(n600) );
  XNOR2_X1 U692 ( .A(n601), .B(KEYINPUT77), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n763), .A2(KEYINPUT47), .ZN(n602) );
  XOR2_X1 U694 ( .A(KEYINPUT86), .B(n602), .Z(n614) );
  NAND2_X1 U695 ( .A1(n746), .A2(n603), .ZN(n619) );
  INV_X1 U696 ( .A(n619), .ZN(n604) );
  AND2_X1 U697 ( .A1(n605), .A2(n604), .ZN(n607) );
  INV_X1 U698 ( .A(n733), .ZN(n606) );
  NAND2_X1 U699 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U700 ( .A1(n608), .A2(n621), .ZN(n612) );
  NAND2_X1 U701 ( .A1(n553), .A2(n718), .ZN(n609) );
  XOR2_X1 U702 ( .A(KEYINPUT30), .B(n609), .Z(n611) );
  AND2_X1 U703 ( .A1(n610), .A2(n611), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n612), .A2(n618), .ZN(n656) );
  NAND2_X1 U705 ( .A1(n715), .A2(KEYINPUT47), .ZN(n613) );
  INV_X1 U706 ( .A(n618), .ZN(n624) );
  INV_X1 U707 ( .A(KEYINPUT38), .ZN(n620) );
  XNOR2_X1 U708 ( .A(n621), .B(n620), .ZN(n717) );
  XOR2_X1 U709 ( .A(KEYINPUT92), .B(KEYINPUT39), .Z(n625) );
  XNOR2_X1 U710 ( .A(n626), .B(n625), .ZN(n642) );
  INV_X1 U711 ( .A(n627), .ZN(n768) );
  NAND2_X1 U712 ( .A1(n642), .A2(n768), .ZN(n629) );
  INV_X1 U713 ( .A(KEYINPUT42), .ZN(n633) );
  INV_X1 U714 ( .A(KEYINPUT113), .ZN(n630) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n637), .A2(n552), .ZN(n639) );
  XOR2_X1 U717 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n638) );
  XNOR2_X1 U718 ( .A(n639), .B(n638), .ZN(n641) );
  INV_X1 U719 ( .A(n621), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n658) );
  AND2_X1 U721 ( .A1(n642), .A2(n770), .ZN(n775) );
  NOR2_X1 U722 ( .A1(n658), .A2(n775), .ZN(n643) );
  INV_X1 U723 ( .A(KEYINPUT89), .ZN(n644) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n647), .A2(KEYINPUT2), .ZN(n648) );
  BUF_X2 U726 ( .A(n649), .Z(n782) );
  INV_X1 U727 ( .A(n650), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n651), .A2(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n696), .A2(G478), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(G143), .ZN(G45) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(G42) );
  XNOR2_X1 U733 ( .A(n659), .B(G101), .ZN(G3) );
  XNOR2_X1 U734 ( .A(n660), .B(G119), .ZN(G21) );
  XNOR2_X1 U735 ( .A(KEYINPUT127), .B(KEYINPUT126), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n661), .B(n670), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n670), .B(G227), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n671), .A2(G900), .ZN(n672) );
  NAND2_X1 U743 ( .A1(G953), .A2(n672), .ZN(n673) );
  NAND2_X1 U744 ( .A1(n674), .A2(n673), .ZN(G72) );
  XOR2_X1 U745 ( .A(n676), .B(G137), .Z(G39) );
  XNOR2_X1 U746 ( .A(G110), .B(KEYINPUT116), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n379), .B(n677), .ZN(G12) );
  XNOR2_X1 U748 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(KEYINPUT55), .ZN(n680) );
  XNOR2_X1 U750 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U753 ( .A(KEYINPUT115), .B(KEYINPUT62), .ZN(n686) );
  XNOR2_X1 U754 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U756 ( .A(KEYINPUT93), .B(KEYINPUT63), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n692), .B(n691), .ZN(G57) );
  XOR2_X1 U758 ( .A(n693), .B(G122), .Z(G24) );
  NOR2_X1 U759 ( .A1(n695), .A2(n701), .ZN(G66) );
  NAND2_X1 U760 ( .A1(n696), .A2(G469), .ZN(n700) );
  XOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  XNOR2_X1 U762 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U763 ( .A(n700), .B(n699), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(G54) );
  NOR2_X1 U765 ( .A1(n381), .A2(KEYINPUT2), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n704), .A2(KEYINPUT87), .ZN(n709) );
  INV_X1 U767 ( .A(KEYINPUT87), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n705), .A2(KEYINPUT2), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n661), .A2(n706), .ZN(n707) );
  NOR2_X1 U770 ( .A1(n782), .A2(n707), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U773 ( .A(n712), .B(KEYINPUT88), .ZN(n755) );
  BUF_X1 U774 ( .A(n713), .Z(n714) );
  NOR2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n723) );
  INV_X1 U776 ( .A(n717), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n719), .A2(n718), .ZN(n721) );
  NOR2_X1 U778 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U780 ( .A(KEYINPUT119), .B(n724), .Z(n725) );
  NOR2_X1 U781 ( .A1(n714), .A2(n725), .ZN(n726) );
  XNOR2_X1 U782 ( .A(n726), .B(KEYINPUT120), .ZN(n744) );
  XOR2_X1 U783 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n731) );
  INV_X1 U784 ( .A(n727), .ZN(n728) );
  NAND2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n732), .A2(n553), .ZN(n736) );
  NAND2_X1 U788 ( .A1(n382), .A2(n733), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n734), .B(KEYINPUT50), .ZN(n735) );
  NAND2_X1 U790 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U791 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U792 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(n742) );
  INV_X1 U794 ( .A(n750), .ZN(n741) );
  NOR2_X1 U795 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U797 ( .A(n745), .B(KEYINPUT52), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n746), .A2(G952), .ZN(n747) );
  NOR2_X1 U799 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U800 ( .A1(n749), .A2(G953), .ZN(n753) );
  INV_X1 U801 ( .A(n714), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U804 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n756) );
  XNOR2_X1 U805 ( .A(n757), .B(n756), .ZN(G75) );
  NAND2_X1 U806 ( .A1(n759), .A2(n768), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(G104), .ZN(G6) );
  XOR2_X1 U808 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n761) );
  NAND2_X1 U809 ( .A1(n759), .A2(n770), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U811 ( .A(G107), .B(n762), .ZN(G9) );
  XOR2_X1 U812 ( .A(G128), .B(KEYINPUT29), .Z(n765) );
  INV_X1 U813 ( .A(n763), .ZN(n766) );
  NAND2_X1 U814 ( .A1(n766), .A2(n770), .ZN(n764) );
  XNOR2_X1 U815 ( .A(n765), .B(n764), .ZN(G30) );
  NAND2_X1 U816 ( .A1(n766), .A2(n768), .ZN(n767) );
  XNOR2_X1 U817 ( .A(n767), .B(G146), .ZN(G48) );
  NAND2_X1 U818 ( .A1(n771), .A2(n768), .ZN(n769) );
  XNOR2_X1 U819 ( .A(n769), .B(G113), .ZN(G15) );
  NAND2_X1 U820 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U821 ( .A(n772), .B(G116), .ZN(G18) );
  XNOR2_X1 U822 ( .A(n773), .B(G125), .ZN(n774) );
  XNOR2_X1 U823 ( .A(n774), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U824 ( .A(G134), .B(n775), .Z(G36) );
  XNOR2_X1 U825 ( .A(n776), .B(G101), .ZN(n777) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(n781) );
  NAND2_X1 U827 ( .A1(n779), .A2(G953), .ZN(n780) );
  AND2_X1 U828 ( .A1(n781), .A2(n780), .ZN(n793) );
  INV_X1 U829 ( .A(n782), .ZN(n784) );
  NAND2_X1 U830 ( .A1(n784), .A2(n783), .ZN(n790) );
  XOR2_X1 U831 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n786) );
  NAND2_X1 U832 ( .A1(G224), .A2(G953), .ZN(n785) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(n787) );
  NAND2_X1 U834 ( .A1(G898), .A2(n787), .ZN(n788) );
  XNOR2_X1 U835 ( .A(n788), .B(KEYINPUT124), .ZN(n789) );
  NAND2_X1 U836 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U837 ( .A(n791), .B(KEYINPUT125), .Z(n792) );
  XNOR2_X1 U838 ( .A(n793), .B(n792), .ZN(G69) );
  XOR2_X1 U839 ( .A(G131), .B(n794), .Z(G33) );
endmodule

