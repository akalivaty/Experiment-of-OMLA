//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n207), .A2(new_n208), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n214), .B1(new_n208), .B2(new_n207), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0023(.A(G238), .B(G244), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT2), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n228), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G58), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(KEYINPUT6), .ZN(new_n242));
  INV_X1    g0042(.A(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G97), .A2(G107), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n244), .A2(KEYINPUT6), .A3(G97), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n249), .A2(G20), .B1(G77), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT7), .B1(new_n254), .B2(new_n212), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT7), .ZN(new_n256));
  NOR4_X1   g0056(.A1(new_n252), .A2(new_n253), .A3(new_n256), .A4(G20), .ZN(new_n257));
  OAI21_X1  g0057(.A(G107), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n211), .B1(new_n205), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(new_n212), .A3(G1), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(G97), .C1(new_n263), .C2(new_n264), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n243), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT79), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(KEYINPUT79), .A3(new_n272), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT5), .A2(G41), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT5), .A2(G41), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n260), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n279), .A2(new_n281), .A3(G274), .A4(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n277), .B2(new_n278), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  INV_X1    g0086(.A(G257), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(G244), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT4), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n254), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G250), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT4), .A4(G244), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G283), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n295), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n288), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G200), .ZN(new_n304));
  AOI211_X1 g0104(.A(G190), .B(new_n288), .C1(new_n301), .C2(new_n302), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n266), .B(new_n276), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n275), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n266), .B1(new_n307), .B2(new_n273), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n311), .B(new_n288), .C1(new_n301), .C2(new_n302), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n308), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n270), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n265), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT81), .B(G87), .Z(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n246), .ZN(new_n321));
  NAND3_X1  g0121(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n212), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n323), .A2(KEYINPUT80), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(KEYINPUT80), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n260), .A2(new_n243), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT19), .B1(new_n327), .B2(new_n212), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n254), .A2(G20), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(G68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n265), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(new_n268), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n319), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n292), .A2(G244), .A3(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G116), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n291), .A2(new_n292), .ZN(new_n337));
  INV_X1    g0137(.A(G238), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n302), .ZN(new_n340));
  OAI21_X1  g0140(.A(G250), .B1(new_n282), .B2(G1), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n283), .A2(G274), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n302), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n311), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n339), .B2(new_n302), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n309), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n334), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(G200), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n331), .A2(new_n265), .B1(new_n268), .B2(new_n317), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(G190), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n316), .A2(G87), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n350), .A2(new_n351), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT82), .B1(new_n314), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n349), .A2(new_n354), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT82), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n357), .A2(new_n358), .A3(new_n306), .A4(new_n313), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n260), .A2(G97), .ZN(new_n360));
  AOI21_X1  g0160(.A(G20), .B1(new_n360), .B2(new_n300), .ZN(new_n361));
  INV_X1    g0161(.A(G116), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n212), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n261), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT20), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n268), .A2(new_n362), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n263), .A2(new_n264), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n270), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n366), .B(new_n367), .C1(new_n362), .C2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n292), .A2(G264), .A3(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G303), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n372), .B2(new_n292), .C1(new_n337), .C2(new_n287), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n302), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n281), .A2(G274), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n285), .ZN(new_n376));
  INV_X1    g0176(.A(new_n286), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(G270), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n370), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(new_n370), .A3(G179), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n309), .B1(new_n374), .B2(new_n378), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n370), .A2(KEYINPUT21), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT21), .B1(new_n370), .B2(new_n387), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n356), .A2(new_n359), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n212), .A2(G1), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n265), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G50), .ZN(new_n395));
  INV_X1    g0195(.A(G50), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n268), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT8), .B(G58), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n212), .A2(G33), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n401));
  INV_X1    g0201(.A(G150), .ZN(new_n402));
  INV_X1    g0202(.A(new_n250), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n265), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n395), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n406), .A2(KEYINPUT9), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(KEYINPUT9), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT71), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n297), .A2(G223), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G222), .ZN(new_n412));
  INV_X1    g0212(.A(G77), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n337), .A2(new_n412), .B1(new_n413), .B2(new_n292), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT67), .ZN(new_n415));
  OR3_X1    g0215(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n411), .B2(new_n414), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n302), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT65), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(G1), .B1(new_n280), .B2(new_n282), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT65), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n375), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n281), .A2(new_n419), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(G226), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G190), .ZN(new_n429));
  AOI21_X1  g0229(.A(G200), .B1(new_n418), .B2(new_n427), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n409), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT10), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n311), .B2(new_n428), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n406), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT69), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(KEYINPUT69), .A3(new_n406), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n424), .B1(G244), .B2(new_n426), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n337), .A2(new_n227), .B1(new_n244), .B2(new_n292), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(G238), .B2(new_n297), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(new_n281), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G169), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n311), .B2(new_n443), .ZN(new_n445));
  INV_X1    g0245(.A(new_n268), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G77), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n394), .B2(G77), .ZN(new_n448));
  INV_X1    g0248(.A(new_n398), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT70), .ZN(new_n451));
  OR3_X1    g0251(.A1(new_n317), .A2(new_n451), .A3(new_n399), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n317), .B2(new_n399), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n265), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n443), .A2(new_n383), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G190), .B2(new_n443), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n455), .A3(new_n448), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n432), .A2(new_n439), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT73), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n292), .A2(G226), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n327), .B1(new_n463), .B2(new_n291), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n297), .A2(G232), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n302), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT13), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n424), .B1(G238), .B2(new_n426), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n281), .B1(new_n464), .B2(new_n465), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n423), .A2(new_n421), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G274), .A3(new_n281), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n338), .B2(new_n425), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT13), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n462), .B1(new_n476), .B2(new_n311), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n470), .A2(new_n475), .A3(KEYINPUT73), .A4(G179), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT14), .B1(new_n476), .B2(G169), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(KEYINPUT14), .A3(G169), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G68), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n413), .B2(new_n399), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n265), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(KEYINPUT11), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(KEYINPUT11), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n267), .A2(G1), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G20), .A3(new_n484), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT12), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n394), .A2(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT72), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n483), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n470), .A2(new_n475), .A3(new_n381), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n476), .A2(new_n383), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n461), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT16), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n256), .B1(new_n292), .B2(G20), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n484), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G58), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n484), .ZN(new_n509));
  OAI21_X1  g0309(.A(G20), .B1(new_n509), .B2(new_n201), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n250), .A2(G159), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n504), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(G68), .B1(new_n255), .B2(new_n257), .ZN(new_n514));
  INV_X1    g0314(.A(new_n512), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(KEYINPUT16), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n516), .A3(new_n265), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n446), .A2(new_n398), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n394), .B2(new_n398), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n292), .A2(G226), .A3(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G87), .ZN(new_n523));
  INV_X1    g0323(.A(G223), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n337), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n302), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n426), .A2(G232), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n473), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n383), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n425), .A2(new_n227), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT75), .B1(new_n424), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT75), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n473), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n531), .A2(new_n533), .A3(new_n381), .A4(new_n526), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n521), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n521), .A2(new_n535), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n517), .A2(KEYINPUT74), .A3(new_n519), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT74), .B1(new_n517), .B2(new_n519), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n528), .A2(new_n309), .ZN(new_n546));
  AOI21_X1  g0346(.A(G179), .B1(new_n525), .B2(new_n302), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n531), .A3(new_n533), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT76), .B1(new_n550), .B2(KEYINPUT18), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(KEYINPUT76), .A3(KEYINPUT18), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT78), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n555), .A2(KEYINPUT78), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n503), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n490), .A2(G20), .A3(new_n244), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n559), .B2(new_n560), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n369), .B2(new_n244), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n212), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n244), .A2(KEYINPUT23), .A3(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n329), .A2(new_n573), .A3(G87), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n292), .A2(new_n212), .A3(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT22), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n577), .A2(KEYINPUT24), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n368), .B1(new_n577), .B2(KEYINPUT24), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n566), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G257), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT84), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n292), .A2(new_n584), .A3(G257), .A4(G1698), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n291), .A2(new_n292), .A3(G250), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n302), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n285), .A2(G264), .A3(new_n281), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n311), .A3(new_n591), .A4(new_n284), .ZN(new_n592));
  AOI211_X1 g0392(.A(new_n590), .B(new_n376), .C1(new_n588), .C2(new_n302), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(KEYINPUT85), .C1(new_n593), .C2(G169), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n589), .A2(new_n591), .A3(new_n284), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n309), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT85), .B1(new_n597), .B2(new_n592), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n581), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT86), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT87), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT85), .ZN(new_n603));
  INV_X1    g0403(.A(new_n592), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n590), .B1(new_n588), .B2(new_n302), .ZN(new_n605));
  AOI21_X1  g0405(.A(G169), .B1(new_n605), .B2(new_n284), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n594), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(KEYINPUT86), .A3(new_n581), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n593), .A2(G200), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n596), .A2(G190), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n580), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n601), .A2(new_n602), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n601), .A2(new_n609), .A3(new_n612), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT87), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n392), .B(new_n558), .C1(new_n613), .C2(new_n615), .ZN(G372));
  AND2_X1   g0416(.A1(new_n531), .A2(new_n533), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(new_n547), .B1(new_n309), .B2(new_n528), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n520), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT18), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT18), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n621), .A3(new_n520), .ZN(new_n622));
  INV_X1    g0422(.A(new_n497), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n501), .A2(new_n500), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n457), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n499), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n620), .B(new_n622), .C1(new_n627), .C2(new_n543), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n432), .B1(new_n437), .B2(new_n438), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n303), .A2(G179), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n309), .B2(new_n303), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n349), .A3(new_n308), .A4(new_n354), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT89), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n313), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n357), .A2(new_n635), .A3(new_n636), .A4(KEYINPUT26), .ZN(new_n637));
  OR3_X1    g0437(.A1(new_n347), .A2(KEYINPUT88), .A3(new_n383), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT88), .B1(new_n347), .B2(new_n383), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n349), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n313), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n634), .B(new_n637), .C1(KEYINPUT26), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n349), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n389), .A2(new_n390), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n581), .A2(new_n592), .A3(new_n597), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n351), .A2(new_n353), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n352), .A3(new_n639), .A4(new_n638), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n612), .A2(new_n650), .A3(new_n306), .A4(new_n313), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n645), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n629), .B1(new_n558), .B2(new_n653), .ZN(G369));
  NAND2_X1  g0454(.A1(new_n490), .A2(new_n212), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT27), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT90), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n656), .A2(KEYINPUT90), .A3(new_n657), .ZN(new_n660));
  OAI221_X1 g0460(.A(G213), .B1(KEYINPUT27), .B2(new_n655), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n581), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT91), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n615), .B2(new_n613), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n599), .A2(new_n663), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n370), .ZN(new_n670));
  INV_X1    g0470(.A(new_n646), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n385), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n646), .A2(new_n370), .A3(new_n664), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n647), .A2(new_n664), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n646), .A2(new_n664), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n667), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n206), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G1), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n320), .A2(new_n362), .A3(new_n246), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n209), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n642), .A2(new_n633), .A3(new_n313), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT94), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n633), .B2(new_n632), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT94), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n645), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT86), .B1(new_n608), .B2(new_n581), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n600), .B(new_n580), .C1(new_n607), .C2(new_n594), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n646), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n651), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n664), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n664), .B1(new_n644), .B2(new_n652), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(KEYINPUT29), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n615), .A2(new_n613), .ZN(new_n706));
  INV_X1    g0506(.A(new_n392), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n663), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n380), .A2(G179), .A3(new_n347), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n301), .A2(new_n302), .ZN(new_n710));
  INV_X1    g0510(.A(new_n288), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n712), .A2(KEYINPUT93), .A3(new_n596), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT93), .B1(new_n712), .B2(new_n596), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT92), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n605), .A2(new_n717), .A3(new_n347), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n380), .A2(new_n718), .A3(G179), .A4(new_n303), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n605), .B2(new_n347), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n712), .A2(new_n311), .A3(new_n379), .ZN(new_n722));
  INV_X1    g0522(.A(new_n720), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n723), .A4(new_n718), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n715), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n664), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n675), .B1(new_n708), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n705), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n690), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(new_n267), .A2(G20), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G45), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n686), .A2(G1), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT96), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n211), .B1(G20), .B2(new_n309), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n210), .A2(G45), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n237), .B2(G45), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n684), .A2(new_n292), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n684), .A2(new_n254), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G355), .B1(new_n362), .B2(new_n684), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n747), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n381), .A2(G20), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n311), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n383), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT99), .Z(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(G311), .B1(new_n768), .B2(G283), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G179), .A2(G200), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n212), .B1(new_n770), .B2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n212), .A2(new_n381), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n311), .A2(new_n383), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G326), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n254), .B1(new_n771), .B2(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n766), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n773), .A2(new_n759), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n372), .A2(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n758), .A2(new_n770), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n777), .B(new_n781), .C1(G329), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n758), .A2(new_n774), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n785), .A2(new_n786), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT33), .B(G317), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT101), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n769), .B(new_n784), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n790), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n794), .A2(G68), .B1(new_n768), .B2(G107), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n320), .A2(new_n778), .B1(new_n779), .B2(new_n508), .ZN(new_n796));
  INV_X1    g0596(.A(new_n775), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n254), .B(new_n796), .C1(G50), .C2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n795), .B(new_n798), .C1(new_n413), .C2(new_n764), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n801));
  OR3_X1    g0601(.A1(new_n782), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n782), .B2(new_n800), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n243), .C2(new_n771), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n793), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n741), .B(new_n756), .C1(new_n805), .C2(new_n745), .ZN(new_n806));
  INV_X1    g0606(.A(new_n674), .ZN(new_n807));
  INV_X1    g0607(.A(new_n744), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n741), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n807), .A2(G330), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT95), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n811), .B1(new_n812), .B2(new_n677), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(G396));
  INV_X1    g0616(.A(new_n745), .ZN(new_n817));
  INV_X1    g0617(.A(new_n779), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G137), .A2(new_n797), .B1(new_n818), .B2(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n819), .B1(new_n790), .B2(new_n402), .C1(new_n800), .C2(new_n764), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n768), .A2(G68), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n396), .B2(new_n778), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT103), .ZN(new_n824));
  INV_X1    g0624(.A(new_n771), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G58), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n254), .B1(new_n783), .B2(G132), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n244), .A2(new_n778), .B1(new_n779), .B2(new_n772), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n254), .B1(new_n771), .B2(new_n243), .C1(new_n782), .C2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(G303), .C2(new_n797), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n765), .A2(G116), .B1(new_n768), .B2(G87), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n832), .B(new_n833), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n828), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n817), .B1(new_n840), .B2(KEYINPUT104), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(KEYINPUT104), .B2(new_n840), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n745), .A2(new_n742), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n842), .B(new_n810), .C1(G77), .C2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n456), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n460), .B1(new_n846), .B2(new_n663), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n457), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n445), .A2(new_n456), .A3(new_n663), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(new_n742), .B2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT105), .Z(new_n852));
  XNOR2_X1  g0652(.A(new_n704), .B(new_n850), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(new_n731), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n731), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n854), .A2(new_n855), .A3(new_n810), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n736), .A2(new_n269), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n497), .B(new_n664), .C1(new_n483), .C2(new_n502), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n497), .A2(new_n664), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n476), .A2(G169), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT14), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n481), .B1(new_n477), .B2(new_n478), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n625), .B(new_n861), .C1(new_n865), .C2(new_n623), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n850), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT31), .B1(new_n725), .B2(new_n664), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n729), .B1(new_n870), .B2(KEYINPUT110), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT110), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n872), .B(KEYINPUT31), .C1(new_n725), .C2(new_n664), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n869), .B1(new_n708), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT40), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n536), .A2(new_n619), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n520), .A2(new_n662), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT74), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n520), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n517), .A2(KEYINPUT74), .A3(new_n519), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n618), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n662), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n536), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n888), .C1(new_n555), .C2(new_n878), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n544), .A2(new_n545), .A3(new_n661), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n877), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT109), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n887), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n620), .A2(new_n622), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n891), .B1(new_n543), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n892), .B2(new_n887), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n890), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n876), .B1(new_n889), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n875), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT76), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n884), .B2(new_n621), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n884), .A2(new_n621), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n554), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n543), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n878), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n888), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n890), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n889), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n889), .B2(new_n909), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n875), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n901), .B1(new_n913), .B2(new_n876), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n392), .B(new_n664), .C1(new_n615), .C2(new_n613), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n728), .A2(new_n872), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n870), .A2(KEYINPUT110), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n729), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n558), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n914), .B(new_n920), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(G330), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT111), .Z(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n849), .B(KEYINPUT106), .Z(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n704), .B2(new_n868), .ZN(new_n926));
  INV_X1    g0726(.A(new_n867), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n911), .B2(new_n912), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n498), .A2(new_n664), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT108), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n889), .A2(new_n933), .A3(new_n899), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n889), .B2(new_n909), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n895), .A2(new_n661), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n929), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n629), .B1(new_n705), .B2(new_n558), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n859), .B1(new_n924), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n924), .B2(new_n940), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n209), .A2(new_n413), .A3(new_n509), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n484), .A2(G50), .ZN(new_n944));
  OAI211_X1 g0744(.A(G1), .B(new_n267), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(G116), .B(new_n213), .C1(new_n249), .C2(KEYINPUT35), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(KEYINPUT35), .B2(new_n249), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT36), .Z(new_n948));
  NAND3_X1  g0748(.A1(new_n942), .A2(new_n945), .A3(new_n948), .ZN(G367));
  INV_X1    g0749(.A(KEYINPUT113), .ZN(new_n950));
  INV_X1    g0750(.A(new_n669), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n664), .A2(new_n308), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n306), .A2(new_n313), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n313), .B2(new_n663), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(new_n681), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT42), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(KEYINPUT42), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n313), .B1(new_n699), .B2(new_n953), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n663), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n950), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n950), .A3(new_n962), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n663), .A2(new_n649), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n645), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n642), .C2(new_n967), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n966), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n971), .B(KEYINPUT43), .Z(new_n974));
  NAND3_X1  g0774(.A1(new_n964), .A2(new_n965), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n678), .A2(new_n954), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n685), .B(KEYINPUT41), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n667), .A2(new_n681), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n951), .B2(new_n681), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n676), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n734), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n682), .A2(new_n954), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n682), .A2(new_n954), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n679), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n990), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n678), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n985), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n980), .B1(new_n994), .B2(new_n734), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n737), .A2(G1), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n978), .B(new_n979), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n778), .A2(new_n362), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  INV_X1    g0799(.A(new_n837), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(G294), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT114), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n254), .B1(new_n771), .B2(new_n244), .C1(new_n767), .C2(new_n243), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n783), .A2(G317), .B1(new_n818), .B2(G303), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n830), .B2(new_n775), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G283), .C2(new_n765), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1011));
  INV_X1    g0811(.A(G137), .ZN(new_n1012));
  INV_X1    g0812(.A(G143), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n782), .A2(new_n1012), .B1(new_n775), .B2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n767), .A2(new_n413), .B1(new_n778), .B2(new_n508), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n292), .B1(new_n779), .B2(new_n402), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n771), .A2(new_n484), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n396), .B2(new_n764), .C1(new_n837), .C2(new_n800), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT116), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1010), .A2(new_n1011), .A3(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT117), .Z(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT47), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT47), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n745), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n232), .A2(new_n750), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n747), .B1(new_n684), .B2(new_n318), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n741), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1025), .B(new_n1028), .C1(new_n808), .C2(new_n971), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n997), .A2(new_n1029), .ZN(G387));
  NOR2_X1   g0830(.A1(new_n985), .A2(new_n686), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n734), .B2(new_n983), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n983), .A2(new_n996), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n751), .B1(new_n228), .B2(G45), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n688), .B2(new_n754), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n449), .A2(new_n396), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n282), .B1(new_n484), .B2(new_n413), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1037), .A2(new_n688), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1035), .A2(new_n1039), .B1(G107), .B2(new_n206), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n741), .B1(new_n1040), .B2(new_n746), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n782), .A2(new_n402), .B1(new_n775), .B2(new_n800), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G50), .B2(new_n818), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n778), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n254), .B1(new_n1044), .B2(G77), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(new_n317), .C2(new_n771), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n484), .A2(new_n764), .B1(new_n790), .B2(new_n398), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT118), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(G97), .C2(new_n768), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(KEYINPUT119), .B(G322), .ZN(new_n1050));
  INV_X1    g0850(.A(G317), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n775), .A2(new_n1050), .B1(new_n779), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n765), .B2(G303), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n837), .B2(new_n830), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n778), .A2(new_n772), .B1(new_n771), .B2(new_n838), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT49), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n254), .B1(new_n782), .B2(new_n776), .C1(new_n362), .C2(new_n767), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n1059), .B2(KEYINPUT49), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1049), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1041), .B1(new_n817), .B2(new_n1063), .C1(new_n951), .C2(new_n808), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1032), .A2(new_n1033), .A3(new_n1064), .ZN(G393));
  AND2_X1   g0865(.A1(new_n994), .A2(new_n685), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n993), .A2(new_n991), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n984), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n240), .A2(new_n751), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n746), .B1(new_n243), .B2(new_n206), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n810), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n837), .A2(new_n396), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G150), .A2(new_n797), .B1(new_n818), .B2(G159), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n449), .B2(new_n765), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n292), .B1(new_n778), .B2(new_n484), .C1(new_n782), .C2(new_n1013), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G77), .B2(new_n825), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n768), .A2(G87), .B1(KEYINPUT51), .B2(new_n1074), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n837), .A2(new_n372), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n765), .A2(G294), .B1(new_n768), .B2(G107), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n778), .A2(new_n838), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n254), .B1(new_n782), .B2(new_n1050), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(G116), .C2(new_n825), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n775), .A2(new_n1051), .B1(new_n779), .B2(new_n830), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1073), .A2(new_n1080), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1072), .B1(new_n1089), .B2(new_n745), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n954), .B2(new_n808), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n996), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1067), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1069), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G390));
  NAND2_X1  g0895(.A1(new_n905), .A2(new_n906), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n879), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT38), .B1(new_n1097), .B2(new_n888), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n907), .A2(new_n908), .A3(new_n890), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n889), .A2(new_n899), .A3(new_n933), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n742), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n810), .B1(new_n449), .B2(new_n844), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n837), .A2(new_n244), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n782), .A2(new_n772), .B1(new_n779), .B2(new_n362), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n254), .B1(new_n771), .B2(new_n413), .C1(new_n775), .C2(new_n838), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G87), .C2(new_n1044), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1107), .B(new_n822), .C1(new_n243), .C2(new_n764), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n837), .A2(new_n1012), .ZN(new_n1109));
  INV_X1    g0909(.A(G128), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n767), .A2(new_n396), .B1(new_n775), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n292), .B1(new_n771), .B2(new_n800), .C1(new_n782), .C2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(G132), .C2(new_n818), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n778), .A2(new_n402), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1114), .B(new_n1117), .C1(new_n764), .C2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1104), .A2(new_n1108), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1120), .B2(new_n745), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1102), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n889), .A2(new_n899), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n849), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n702), .B2(new_n848), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1124), .B(new_n931), .C1(new_n1126), .C2(new_n927), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1100), .B(new_n1101), .C1(new_n928), .C2(new_n932), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n868), .A2(G330), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n919), .A2(new_n927), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n850), .B1(new_n866), .B2(new_n860), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n731), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1123), .B1(new_n1136), .B2(new_n1092), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n939), .B1(G330), .B2(new_n920), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n867), .B1(new_n731), .B2(new_n868), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n704), .A2(new_n868), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1131), .A2(new_n1139), .B1(new_n1140), .B2(new_n925), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n927), .B1(new_n919), .B2(new_n1130), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1126), .A3(new_n1134), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(new_n1136), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n686), .B1(new_n1145), .B2(new_n1136), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1137), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  NAND2_X1  g0949(.A1(new_n432), .A2(new_n435), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n662), .A2(new_n406), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT124), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1152), .B(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT125), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n929), .A2(new_n936), .A3(new_n937), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n875), .A2(new_n900), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1133), .B1(new_n915), .B2(new_n918), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT107), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n889), .A2(new_n909), .A3(new_n910), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(G330), .B(new_n1159), .C1(new_n1163), .C2(KEYINPUT40), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n938), .B1(new_n914), .B2(G330), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1157), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n914), .A2(new_n938), .A3(G330), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1157), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n996), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1155), .A2(new_n742), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n741), .B1(new_n396), .B2(new_n843), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n317), .A2(new_n764), .B1(new_n790), .B2(new_n243), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT123), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n254), .A2(new_n280), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n767), .A2(new_n508), .B1(new_n782), .B2(new_n838), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(G77), .C2(new_n1044), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT122), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n775), .A2(new_n362), .B1(new_n779), .B2(new_n244), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1177), .A2(new_n1181), .A3(new_n1017), .A4(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT58), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n818), .A2(G128), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n778), .B2(new_n1118), .C1(new_n1112), .C2(new_n775), .ZN(new_n1186));
  INV_X1    g0986(.A(G132), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1012), .A2(new_n764), .B1(new_n790), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G150), .C2(new_n825), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n260), .B(new_n280), .C1(new_n767), .C2(new_n800), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G124), .B2(new_n783), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1178), .B(new_n396), .C1(G33), .C2(G41), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1183), .A2(KEYINPUT58), .ZN(new_n1197));
  AND4_X1   g0997(.A1(new_n1184), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1174), .B(new_n1175), .C1(new_n817), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1173), .A2(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1138), .B1(new_n1136), .B2(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1170), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT57), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1172), .A2(new_n1207), .A3(new_n1202), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1200), .B1(new_n1209), .B2(new_n685), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(G375));
  OR2_X1    g1011(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n980), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1145), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n927), .A2(new_n742), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n810), .B1(G68), .B2(new_n844), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n292), .B1(new_n771), .B2(new_n396), .C1(new_n767), .C2(new_n508), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1012), .A2(new_n779), .B1(new_n778), .B2(new_n800), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n782), .A2(new_n1110), .B1(new_n775), .B2(new_n1187), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n402), .B2(new_n764), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n837), .A2(new_n1118), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n837), .A2(new_n362), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n765), .A2(G107), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n243), .A2(new_n778), .B1(new_n779), .B2(new_n838), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G303), .B2(new_n783), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n254), .B1(new_n775), .B2(new_n772), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n318), .B2(new_n825), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n768), .A2(G77), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1224), .A2(new_n1226), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1221), .A2(new_n1222), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1216), .B1(new_n1231), .B2(new_n745), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1144), .A2(new_n996), .B1(new_n1215), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1214), .A2(new_n1233), .ZN(G381));
  NOR2_X1   g1034(.A1(G375), .A2(G378), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n997), .A2(new_n1094), .A3(new_n1029), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(G393), .A2(G381), .A3(G384), .A4(G396), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .ZN(G407));
  INV_X1    g1039(.A(G213), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(G343), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1235), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(G409));
  INV_X1    g1043(.A(new_n1200), .ZN(new_n1244));
  OR3_X1    g1044(.A1(new_n1205), .A2(KEYINPUT127), .A3(new_n980), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT127), .B1(new_n1205), .B2(new_n980), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1148), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1210), .B2(G378), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n686), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1251), .A2(KEYINPUT126), .A3(new_n1200), .A4(new_n1148), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1248), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1241), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1233), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1212), .B(KEYINPUT60), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n686), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(G384), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n857), .B(new_n1255), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1253), .A2(new_n1254), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1259), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1260), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1241), .A2(G2897), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G2897), .B(new_n1241), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1209), .A2(new_n685), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(G378), .A3(new_n1244), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1210), .A2(new_n1249), .A3(G378), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1273), .A2(new_n1274), .B1(new_n1148), .B2(new_n1247), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1270), .B1(new_n1275), .B2(new_n1241), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1253), .A2(new_n1277), .A3(new_n1254), .A4(new_n1261), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1263), .A2(new_n1264), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1094), .B1(new_n997), .B2(new_n1029), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(G393), .B(G396), .Z(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1236), .A3(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1237), .B2(new_n1280), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1279), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1254), .B2(new_n1253), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1262), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1262), .A2(new_n1290), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1286), .A2(KEYINPUT61), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1287), .A2(new_n1294), .ZN(G405));
  AND3_X1   g1095(.A1(new_n1284), .A2(new_n1285), .A3(new_n1261), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1261), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1273), .A2(new_n1274), .B1(new_n1148), .B2(G375), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1298), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(G402));
endmodule


