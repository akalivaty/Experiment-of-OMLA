//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n226), .A2(new_n227), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n215), .B1(new_n218), .B2(new_n220), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G58), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n222), .ZN(new_n252));
  OAI21_X1  g0052(.A(G20), .B1(new_n252), .B2(new_n201), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G159), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT72), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT72), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT3), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(new_n210), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n264), .B2(KEYINPUT7), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT72), .B(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(new_n269), .B2(new_n210), .ZN(new_n270));
  OAI211_X1 g0070(.A(KEYINPUT16), .B(new_n257), .C1(new_n265), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n216), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  AOI21_X1  g0074(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n275), .A2(KEYINPUT7), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n262), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT72), .A2(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n261), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n263), .A2(new_n275), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n266), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n222), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n274), .B1(new_n284), .B2(new_n256), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n271), .A2(new_n273), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n251), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n292), .A2(new_n210), .A3(G1), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n273), .B1(new_n209), .B2(G20), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n291), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n286), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G226), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1698), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G223), .B2(G1698), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n263), .B2(new_n260), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n300), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  OAI211_X1 g0108(.A(G1), .B(G13), .C1(new_n262), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G45), .ZN(new_n310));
  AOI21_X1  g0110(.A(G1), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(G274), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(G232), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n307), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G223), .A2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n301), .B2(G1698), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n261), .B1(new_n278), .B2(new_n279), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n267), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n309), .B1(new_n319), .B2(new_n305), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G179), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT73), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT73), .B1(new_n312), .B2(new_n314), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n299), .A2(new_n315), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n298), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT18), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n298), .A2(new_n329), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT75), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n312), .A2(new_n314), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n320), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n307), .A2(new_n337), .A3(new_n338), .A4(new_n322), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n335), .B1(new_n339), .B2(KEYINPUT74), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT74), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n320), .A2(G190), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n325), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n286), .B(new_n297), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n286), .A2(new_n297), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n341), .A3(new_n325), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n339), .A2(KEYINPUT74), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n335), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT17), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n332), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n344), .A2(new_n345), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n350), .A3(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT75), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n331), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(KEYINPUT3), .A2(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n263), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G1698), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G222), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G223), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n360), .B1(new_n224), .B2(new_n358), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n300), .ZN(new_n364));
  INV_X1    g0164(.A(new_n312), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n300), .A2(new_n311), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(G226), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G200), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n338), .B2(new_n368), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT67), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n296), .A2(G50), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G50), .B2(new_n294), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n254), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n210), .A2(G33), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n291), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n273), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT10), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n372), .A2(KEYINPUT10), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n372), .A2(KEYINPUT10), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n378), .B(KEYINPUT9), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n370), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n299), .B2(new_n368), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G179), .B2(new_n368), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G20), .A2(G77), .ZN(new_n390));
  INV_X1    g0190(.A(new_n254), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n390), .B1(new_n287), .B2(new_n391), .C1(new_n376), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n273), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n296), .A2(G77), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(new_n395), .C1(G77), .C2(new_n294), .ZN(new_n396));
  INV_X1    g0196(.A(G232), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n263), .B2(new_n357), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n359), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(new_n206), .B2(new_n358), .C1(new_n361), .C2(new_n223), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n300), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n365), .B1(G244), .B2(new_n366), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n403), .B2(G190), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n333), .B2(new_n403), .ZN(new_n405));
  INV_X1    g0205(.A(G179), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n396), .B1(new_n403), .B2(G169), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n356), .A2(new_n389), .A3(new_n405), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n293), .A2(new_n222), .ZN(new_n412));
  XOR2_X1   g0212(.A(new_n412), .B(KEYINPUT12), .Z(new_n413));
  OAI22_X1  g0213(.A1(new_n391), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n376), .A2(new_n224), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n273), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT11), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n296), .A2(G68), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n413), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  XOR2_X1   g0221(.A(new_n421), .B(KEYINPUT71), .Z(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n365), .B1(G238), .B2(new_n366), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n398), .A2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT68), .ZN(new_n429));
  AOI21_X1  g0229(.A(G1698), .B1(new_n263), .B2(new_n357), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(G226), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n429), .A3(G226), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n300), .B1(new_n434), .B2(KEYINPUT69), .ZN(new_n435));
  INV_X1    g0235(.A(new_n433), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n426), .B(new_n427), .C1(new_n436), .C2(new_n431), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT69), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n424), .B(new_n425), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n434), .A2(KEYINPUT69), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n300), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n424), .B1(new_n444), .B2(new_n425), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n423), .B(G169), .C1(new_n441), .C2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n425), .B1(new_n435), .B2(new_n439), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT13), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(G179), .A3(new_n440), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n440), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n423), .B1(new_n451), .B2(G169), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n422), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(G190), .A3(new_n440), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT70), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n451), .B2(G200), .ZN(new_n456));
  AOI211_X1 g0256(.A(KEYINPUT70), .B(new_n333), .C1(new_n448), .C2(new_n440), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n421), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n411), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(G1698), .B1(new_n260), .B2(new_n263), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(KEYINPUT81), .A3(G257), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n260), .A2(new_n263), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G264), .A2(G1698), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT82), .B(new_n465), .C1(new_n260), .C2(new_n263), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n263), .A2(new_n357), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G303), .ZN(new_n471));
  INV_X1    g0271(.A(G257), .ZN(new_n472));
  AOI211_X1 g0272(.A(new_n472), .B(G1698), .C1(new_n260), .C2(new_n263), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n473), .B2(KEYINPUT81), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n300), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT5), .B(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n310), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n300), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G270), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n309), .A2(G274), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n478), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n299), .B1(new_n475), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n273), .C1(new_n210), .C2(G116), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT20), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n294), .A2(G116), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n209), .A2(G33), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n492), .A2(KEYINPUT77), .ZN(new_n493));
  INV_X1    g0293(.A(new_n273), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(KEYINPUT77), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n294), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n490), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT21), .B1(new_n486), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n464), .A2(G257), .A3(new_n359), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(G303), .B2(new_n470), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT82), .B1(new_n269), .B2(new_n465), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n464), .A2(new_n463), .A3(new_n466), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n462), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n484), .B1(new_n508), .B2(new_n300), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n486), .A2(KEYINPUT21), .B1(new_n509), .B2(G179), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT83), .B1(new_n510), .B2(new_n499), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n505), .A2(new_n506), .B1(new_n473), .B2(KEYINPUT81), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n309), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  OAI211_X1 g0313(.A(KEYINPUT21), .B(G169), .C1(new_n513), .C2(new_n484), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n475), .A2(G179), .A3(new_n485), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n500), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n501), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n472), .A2(G1698), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(G250), .B2(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G294), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n258), .A2(new_n259), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n269), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n300), .B1(new_n479), .B2(G264), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n483), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(G179), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n299), .B2(new_n526), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n206), .A2(G20), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n523), .A2(new_n497), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n533), .B2(G20), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G87), .ZN(new_n536));
  OR4_X1    g0336(.A1(KEYINPUT22), .A2(new_n470), .A3(G20), .A4(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n210), .B(G87), .C1(new_n318), .C2(new_n267), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT22), .B1(new_n538), .B2(KEYINPUT84), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  AOI21_X1  g0340(.A(G20), .B1(new_n260), .B2(new_n263), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G87), .ZN(new_n542));
  OAI211_X1 g0342(.A(KEYINPUT85), .B(new_n537), .C1(new_n539), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(KEYINPUT84), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(new_n540), .A3(G87), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT22), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT85), .B1(new_n547), .B2(new_n537), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n535), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n537), .B1(new_n539), .B2(new_n542), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n543), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n535), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n494), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n529), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n292), .A2(G1), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT86), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT25), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n561), .A2(KEYINPUT25), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(KEYINPUT25), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n558), .A2(new_n563), .A3(new_n559), .A4(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n565), .C1(new_n496), .C2(new_n206), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n528), .B1(new_n557), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n555), .B1(new_n554), .B2(new_n535), .ZN(new_n568));
  AOI211_X1 g0368(.A(KEYINPUT24), .B(new_n534), .C1(new_n553), .C2(new_n543), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n273), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n566), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n526), .B2(new_n338), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G200), .B2(new_n526), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n475), .A2(new_n485), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n500), .B1(new_n575), .B2(G200), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n338), .B2(new_n575), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n519), .A2(new_n567), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n293), .A2(KEYINPUT76), .A3(new_n205), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT76), .B1(new_n293), .B2(new_n205), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n496), .A2(new_n205), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n254), .A2(G77), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G97), .A2(G107), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT6), .B1(new_n207), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n276), .A2(new_n280), .B1(new_n282), .B2(new_n266), .ZN(new_n587));
  OAI221_X1 g0387(.A(new_n582), .B1(new_n586), .B2(new_n210), .C1(new_n587), .C2(new_n206), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n581), .B1(new_n588), .B2(new_n273), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n430), .A2(KEYINPUT4), .A3(G244), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n358), .A2(G250), .A3(G1698), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n487), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(new_n359), .C1(new_n318), .C2(new_n267), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(KEYINPUT78), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT78), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n461), .B2(G244), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n300), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n479), .A2(G257), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n483), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(G179), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n589), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n595), .A2(KEYINPUT78), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n461), .A2(new_n597), .A3(G244), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n594), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n309), .B1(new_n607), .B2(new_n593), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n299), .B1(new_n608), .B2(new_n602), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(G200), .B1(new_n608), .B2(new_n602), .ZN(new_n612));
  INV_X1    g0412(.A(new_n602), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n225), .B(G1698), .C1(new_n260), .C2(new_n263), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT4), .B1(new_n614), .B2(new_n597), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n592), .B1(new_n615), .B2(new_n605), .ZN(new_n616));
  OAI211_X1 g0416(.A(G190), .B(new_n613), .C1(new_n616), .C2(new_n309), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(new_n617), .A3(new_n589), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT79), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT79), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n612), .A2(new_n617), .A3(new_n620), .A4(new_n589), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n611), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n223), .A2(new_n359), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n225), .A2(G1698), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n260), .B2(new_n263), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n300), .B1(new_n626), .B2(new_n532), .ZN(new_n627));
  INV_X1    g0427(.A(G250), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n477), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n482), .A2(new_n477), .B1(new_n309), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n210), .B(G68), .C1(new_n318), .C2(new_n267), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT19), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT80), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT80), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT19), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n205), .B2(new_n376), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n536), .A2(new_n205), .A3(new_n206), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n427), .A2(new_n210), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n635), .A4(new_n637), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n633), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n273), .B1(new_n293), .B2(new_n392), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n494), .A2(new_n294), .A3(new_n493), .A4(new_n495), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G87), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n627), .A2(new_n630), .A3(G190), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n632), .A2(new_n644), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  AOI211_X1 g0448(.A(G20), .B(new_n222), .C1(new_n260), .C2(new_n263), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n639), .A2(new_n642), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n273), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n392), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n392), .A2(new_n293), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n631), .A2(new_n299), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n627), .A2(new_n630), .A3(new_n406), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n622), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n460), .A2(new_n578), .A3(new_n660), .ZN(G372));
  AOI21_X1  g0461(.A(new_n333), .B1(new_n627), .B2(new_n630), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n623), .B(new_n624), .C1(new_n318), .C2(new_n267), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n309), .B1(new_n663), .B2(new_n533), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n482), .A2(new_n477), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n629), .A2(new_n309), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n662), .B1(new_n668), .B2(G190), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT87), .B1(new_n644), .B2(new_n646), .ZN(new_n670));
  AND4_X1   g0470(.A1(KEYINPUT87), .A2(new_n651), .A3(new_n654), .A4(new_n646), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n658), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n570), .B2(new_n573), .ZN(new_n674));
  INV_X1    g0474(.A(new_n528), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n570), .B2(new_n571), .ZN(new_n676));
  INV_X1    g0476(.A(new_n501), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n510), .B2(new_n499), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n622), .B(new_n674), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n658), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n659), .A2(KEYINPUT26), .A3(new_n609), .A4(new_n604), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n672), .A2(new_n604), .A3(new_n658), .A4(new_n609), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n681), .A2(KEYINPUT88), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT88), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n611), .A2(new_n685), .A3(KEYINPUT26), .A4(new_n659), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n680), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n460), .B1(new_n679), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n454), .A2(new_n421), .ZN(new_n689));
  OAI21_X1  g0489(.A(G200), .B1(new_n441), .B2(new_n445), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT70), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n451), .A2(new_n455), .A3(G200), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n453), .B1(new_n693), .B2(new_n410), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n352), .A2(new_n355), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n331), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n381), .A2(new_n385), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n387), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n688), .A2(new_n698), .ZN(G369));
  INV_X1    g0499(.A(KEYINPUT90), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n570), .A2(new_n571), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n559), .A2(new_n210), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT89), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT27), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(G213), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G343), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n567), .A3(new_n574), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n676), .A2(new_n710), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n709), .A2(new_n499), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n678), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n517), .B1(new_n516), .B2(new_n500), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT83), .B(new_n499), .C1(new_n514), .C2(new_n515), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n677), .B(new_n577), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n717), .B1(new_n720), .B2(new_n716), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n700), .B1(new_n715), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n722), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT90), .A3(new_n714), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n567), .A2(new_n710), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n567), .A2(new_n574), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n519), .A2(new_n710), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(G399));
  INV_X1    g0531(.A(new_n213), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G41), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n640), .A2(G116), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n220), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n608), .A2(new_n602), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT91), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n475), .A2(new_n741), .A3(G179), .A4(new_n485), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n668), .A2(new_n525), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n739), .A2(new_n740), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(KEYINPUT92), .B(KEYINPUT30), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n600), .A2(KEYINPUT30), .A3(new_n613), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n739), .A2(new_n747), .A3(new_n742), .A4(new_n743), .ZN(new_n748));
  INV_X1    g0548(.A(new_n740), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n668), .A2(G179), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n749), .A2(new_n526), .A3(new_n575), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n710), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(KEYINPUT31), .B(new_n710), .C1(new_n746), .C2(new_n752), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n619), .A2(new_n621), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n757), .A2(new_n659), .A3(new_n610), .A4(new_n709), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n755), .B(new_n756), .C1(new_n578), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n611), .A2(new_n683), .A3(new_n659), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n682), .A2(KEYINPUT26), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(new_n658), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n673), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n622), .A2(new_n574), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n519), .A2(new_n567), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT29), .B1(new_n767), .B2(new_n710), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n710), .B1(new_n679), .B2(new_n687), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT29), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n760), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n738), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(new_n292), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n209), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n733), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n724), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n721), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n778), .B(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n213), .A2(new_n358), .ZN(new_n782));
  INV_X1    g0582(.A(G355), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n783), .B1(G116), .B2(new_n213), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n732), .A2(new_n464), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n220), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(new_n310), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n246), .A2(new_n310), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n216), .B1(G20), .B2(new_n299), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n781), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n210), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n798), .A2(new_n338), .A3(G200), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n536), .A2(new_n799), .B1(new_n800), .B2(new_n206), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n210), .A2(new_n406), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G190), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(G50), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G190), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n802), .A2(G190), .A3(new_n333), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n358), .B1(new_n811), .B2(new_n251), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n802), .A2(new_n806), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G77), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n338), .A2(G179), .A3(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n210), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n802), .A2(new_n338), .A3(G200), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G97), .A2(new_n818), .B1(new_n820), .B2(G68), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n805), .A2(new_n810), .A3(new_n815), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n811), .ZN(new_n823));
  INV_X1    g0623(.A(new_n807), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n823), .A2(G322), .B1(new_n824), .B2(G329), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n470), .C1(new_n826), .C2(new_n813), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT33), .B(G317), .Z(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n819), .A2(new_n828), .B1(new_n800), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n799), .B(KEYINPUT95), .Z(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G294), .A2(new_n818), .B1(new_n804), .B2(G326), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT94), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n822), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n797), .B1(new_n838), .B2(new_n794), .ZN(new_n839));
  INV_X1    g0639(.A(new_n793), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n721), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n780), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  XNOR2_X1  g0643(.A(new_n409), .B(KEYINPUT100), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(new_n405), .A3(new_n709), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n679), .B2(new_n687), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n710), .A2(new_n396), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n844), .A2(new_n405), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n410), .B2(new_n709), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n847), .B1(new_n769), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n778), .B1(new_n851), .B2(new_n760), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n760), .B2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n794), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n358), .B1(new_n833), .B2(G107), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT96), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G116), .A2(new_n814), .B1(new_n824), .B2(G311), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n522), .B2(new_n811), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n817), .A2(new_n205), .B1(new_n819), .B2(new_n829), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n803), .A2(new_n832), .B1(new_n800), .B2(new_n536), .ZN(new_n860));
  OR4_X1    g0660(.A1(new_n856), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n820), .A2(G150), .B1(new_n804), .B2(G137), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT97), .ZN(new_n863));
  INV_X1    g0663(.A(G143), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n864), .B2(new_n811), .C1(new_n808), .C2(new_n813), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT34), .Z(new_n866));
  INV_X1    g0666(.A(G132), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n464), .B1(new_n867), .B2(new_n807), .C1(new_n251), .C2(new_n817), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n834), .A2(new_n202), .B1(new_n222), .B2(new_n800), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(KEYINPUT98), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(KEYINPUT98), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n861), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT99), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n854), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n873), .B2(new_n872), .ZN(new_n875));
  INV_X1    g0675(.A(new_n781), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n794), .A2(new_n791), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n224), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n875), .B(new_n878), .C1(new_n792), .C2(new_n850), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n853), .A2(new_n879), .ZN(G384));
  NOR2_X1   g0680(.A1(new_n775), .A2(new_n209), .ZN(new_n881));
  INV_X1    g0681(.A(G330), .ZN(new_n882));
  INV_X1    g0682(.A(new_n460), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n759), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT101), .ZN(new_n885));
  OAI21_X1  g0685(.A(G169), .B1(new_n441), .B2(new_n445), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT14), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n449), .A3(new_n446), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n422), .B(new_n710), .C1(new_n693), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n422), .A2(new_n710), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n453), .A2(new_n458), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n759), .A2(new_n850), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n298), .A2(new_n708), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n327), .A2(new_n344), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n326), .A2(new_n708), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n265), .A2(new_n270), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT16), .B1(new_n898), .B2(new_n257), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n271), .A2(new_n273), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n297), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n897), .A2(new_n901), .B1(new_n347), .B2(new_n350), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n896), .B1(new_n902), .B2(new_n895), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n708), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n356), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(KEYINPUT38), .B(new_n903), .C1(new_n356), .C2(new_n904), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT40), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n353), .A2(new_n354), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n298), .B(new_n708), .C1(new_n911), .C2(new_n331), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n327), .A2(new_n344), .A3(new_n894), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n896), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n906), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n759), .A2(new_n918), .A3(new_n892), .A4(new_n850), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n910), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n882), .B1(new_n885), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n885), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n844), .A2(new_n710), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n892), .B1(new_n846), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n907), .A2(new_n908), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n888), .A2(new_n422), .A3(new_n709), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n331), .A2(new_n707), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n927), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n460), .B1(new_n768), .B2(new_n771), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n698), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n881), .B1(new_n923), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n923), .ZN(new_n940));
  INV_X1    g0740(.A(new_n586), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(KEYINPUT35), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(KEYINPUT35), .ZN(new_n943));
  NOR4_X1   g0743(.A1(new_n942), .A2(new_n943), .A3(new_n497), .A4(new_n218), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT36), .Z(new_n945));
  OR3_X1    g0745(.A1(new_n220), .A2(new_n224), .A3(new_n252), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n202), .A2(G68), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n292), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n940), .A2(new_n945), .A3(new_n949), .ZN(G367));
  AND2_X1   g0750(.A1(new_n723), .A2(new_n725), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n622), .B1(new_n589), .B2(new_n709), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n611), .A2(new_n710), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n677), .B1(new_n718), .B2(new_n719), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n956), .A2(new_n567), .A3(new_n574), .A4(new_n709), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n955), .A2(KEYINPUT42), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n676), .A2(new_n757), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n709), .B1(new_n959), .B2(new_n611), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT42), .B1(new_n955), .B2(new_n957), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n670), .A2(new_n671), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n963), .A2(new_n658), .A3(new_n709), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n658), .B(new_n672), .C1(new_n963), .C2(new_n709), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT102), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT43), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT102), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(new_n969), .A3(new_n965), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT103), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT103), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n967), .A2(new_n973), .A3(new_n968), .A4(new_n970), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT104), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n951), .A2(new_n954), .A3(new_n962), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n962), .A2(new_n978), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n723), .A2(new_n725), .A3(new_n954), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n975), .B1(new_n972), .B2(new_n974), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n983), .B1(new_n979), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n733), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT105), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n730), .B2(new_n954), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n676), .A2(new_n709), .ZN(new_n991));
  AND4_X1   g0791(.A1(new_n989), .A2(new_n954), .A3(new_n991), .A4(new_n957), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n730), .A2(new_n989), .A3(new_n954), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n957), .A2(new_n991), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT105), .B1(new_n995), .B2(new_n955), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT45), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT44), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n730), .B2(new_n954), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n993), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n951), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n726), .A2(new_n993), .A3(new_n997), .A4(new_n1001), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n956), .A2(new_n709), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n712), .A2(new_n713), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(KEYINPUT106), .A3(new_n957), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n957), .A2(KEYINPUT106), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n1007), .A2(new_n722), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n722), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1009), .A2(new_n772), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1003), .A2(new_n1004), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n987), .B1(new_n1012), .B2(new_n773), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n986), .B1(new_n1013), .B2(new_n777), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n785), .A2(new_n242), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n796), .B1(new_n732), .B2(new_n652), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n876), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n497), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n833), .A2(G116), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(KEYINPUT46), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n800), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n818), .A2(G107), .B1(new_n1021), .B2(G97), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n522), .B2(new_n819), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G283), .A2(new_n814), .B1(new_n824), .B2(G317), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n832), .B2(new_n811), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n269), .B1(new_n826), .B2(new_n803), .ZN(new_n1026));
  NOR4_X1   g0826(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT107), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT107), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n823), .A2(G150), .B1(new_n824), .B2(G137), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1030), .B(new_n358), .C1(new_n202), .C2(new_n813), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n820), .A2(G159), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n251), .B2(new_n799), .C1(new_n222), .C2(new_n817), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n803), .A2(new_n864), .B1(new_n800), .B2(new_n224), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT108), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1028), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT109), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT47), .Z(new_n1039));
  OAI221_X1 g0839(.A(new_n1017), .B1(new_n840), .B2(new_n966), .C1(new_n1039), .C2(new_n854), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1014), .A2(new_n1040), .ZN(G387));
  NOR2_X1   g0841(.A1(new_n239), .A2(new_n310), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n287), .A2(G50), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT50), .Z(new_n1044));
  OAI211_X1 g0844(.A(new_n735), .B(new_n310), .C1(new_n222), .C2(new_n224), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n785), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1042), .B1(KEYINPUT110), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT110), .B2(new_n1046), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(G107), .B2(new_n213), .C1(new_n735), .C2(new_n782), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n795), .ZN(new_n1050));
  INV_X1    g0850(.A(G150), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n813), .A2(new_n222), .B1(new_n807), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G50), .B2(new_n823), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n820), .A2(new_n290), .A3(new_n289), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n269), .B1(G97), .B2(new_n1021), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n652), .A2(new_n818), .B1(new_n804), .B2(G159), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n224), .C2(new_n799), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n464), .B1(G326), .B2(new_n824), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n817), .A2(new_n829), .B1(new_n799), .B2(new_n522), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n823), .A2(G317), .B1(new_n814), .B2(G303), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n804), .A2(G322), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n826), .C2(new_n819), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1059), .B1(new_n497), .B2(new_n800), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1058), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n794), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1050), .A2(new_n1071), .A3(new_n781), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n715), .B2(new_n793), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n777), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1011), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n733), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1074), .A2(new_n773), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  NAND2_X1  g0879(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1076), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n733), .A3(new_n1012), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1003), .A2(new_n777), .A3(new_n1004), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n823), .A2(G311), .B1(new_n804), .B2(G317), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n358), .B1(new_n824), .B2(G322), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n522), .B2(new_n813), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n819), .A2(new_n832), .B1(new_n800), .B2(new_n206), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n817), .A2(new_n497), .B1(new_n799), .B2(new_n829), .ZN(new_n1089));
  OR4_X1    g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n811), .A2(new_n808), .B1(new_n803), .B2(new_n1051), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n813), .A2(new_n287), .B1(new_n807), .B2(new_n864), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n269), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n817), .A2(new_n224), .B1(new_n799), .B2(new_n222), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n819), .A2(new_n202), .B1(new_n800), .B2(new_n536), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n854), .B1(new_n1090), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n786), .A2(new_n249), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n796), .B(new_n1100), .C1(G97), .C2(new_n732), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1099), .A2(new_n876), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n954), .B2(new_n840), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1082), .A2(new_n1104), .ZN(G390));
  NAND4_X1  g0905(.A1(new_n759), .A2(new_n892), .A3(G330), .A4(new_n850), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n925), .A2(KEYINPUT111), .A3(new_n931), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT111), .B1(new_n925), .B2(new_n931), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n929), .A2(new_n930), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n918), .A2(new_n931), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n763), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n956), .A2(new_n676), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n622), .A2(new_n574), .A3(new_n764), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n844), .A2(new_n405), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n709), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n924), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1112), .B1(new_n1120), .B2(new_n892), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1107), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n678), .B1(new_n701), .B2(new_n528), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n687), .B1(new_n1123), .B2(new_n1115), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n845), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n924), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n889), .A2(new_n891), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n931), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT111), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n929), .A2(new_n930), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n925), .A2(KEYINPUT111), .A3(new_n931), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1121), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1106), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1122), .A2(new_n777), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n876), .B1(new_n291), .B2(new_n877), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT113), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n811), .A2(new_n497), .B1(new_n807), .B2(new_n522), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n358), .B(new_n1139), .C1(G97), .C2(new_n814), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n833), .A2(G87), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n818), .A2(G77), .B1(new_n1021), .B2(G68), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n820), .A2(G107), .B1(new_n804), .B2(G283), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n813), .A2(new_n1145), .B1(new_n807), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n470), .B(new_n1147), .C1(G132), .C2(new_n823), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n799), .A2(new_n1051), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G137), .A2(new_n820), .B1(new_n1021), .B2(G50), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G159), .A2(new_n818), .B1(new_n804), .B2(G128), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n854), .B1(new_n1144), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1138), .A2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT114), .Z(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1110), .B2(new_n792), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1136), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1122), .A2(new_n1135), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n760), .A2(new_n460), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n936), .A2(new_n1160), .A3(new_n698), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n755), .A2(new_n756), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n567), .A2(new_n574), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1163), .A2(new_n720), .A3(new_n758), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n850), .C1(new_n1162), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1127), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n765), .A2(new_n766), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n710), .B1(new_n1167), .B2(new_n1113), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n924), .B1(new_n1168), .B2(new_n1117), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1169), .A3(KEYINPUT112), .A4(new_n1106), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(new_n1169), .A3(new_n1106), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT112), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1126), .B1(new_n1166), .B2(new_n1106), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1161), .B(new_n1170), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n734), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1128), .A2(new_n1129), .B1(new_n929), .B2(new_n930), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1107), .B(new_n1121), .C1(new_n1177), .C2(new_n1132), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1106), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1175), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1158), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1161), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT117), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n707), .A2(new_n378), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n388), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT116), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1191), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n381), .A2(new_n385), .A3(new_n387), .A4(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1193), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1190), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1198), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1189), .A3(new_n1196), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1188), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n893), .A2(new_n909), .B1(new_n919), .B2(KEYINPUT40), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n882), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1202), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n921), .A2(G330), .A3(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1204), .A2(new_n1206), .A3(new_n935), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n935), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1185), .B1(new_n1187), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1161), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n927), .A2(new_n933), .A3(new_n934), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1205), .B1(new_n921), .B2(G330), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n882), .B(new_n1202), .C1(new_n910), .C2(new_n920), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1204), .A2(new_n1206), .A3(new_n935), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1185), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n734), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1210), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n777), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n791), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1146), .A2(new_n803), .B1(new_n819), .B2(new_n867), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n823), .A2(G128), .B1(new_n814), .B2(G137), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n799), .B2(new_n1145), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G150), .C2(new_n818), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1021), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n824), .C2(G124), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1021), .A2(G58), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n205), .B2(new_n819), .C1(new_n497), .C2(new_n803), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n823), .A2(G107), .B1(new_n824), .B2(G283), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n392), .B2(new_n813), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n269), .A2(new_n308), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n817), .A2(new_n222), .B1(new_n799), .B2(new_n224), .ZN(new_n1238));
  OR4_X1    g1038(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(KEYINPUT115), .B(KEYINPUT58), .Z(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1237), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1232), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n794), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n777), .B(new_n733), .C1(new_n202), .C2(new_n877), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1222), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1220), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1219), .A2(new_n1250), .ZN(G375));
  OAI21_X1  g1051(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1186), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n987), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1175), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT118), .Z(new_n1256));
  NAND2_X1  g1056(.A1(new_n1127), .A2(new_n791), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n794), .A2(G68), .A3(new_n791), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n811), .A2(new_n829), .B1(new_n807), .B2(new_n832), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n358), .B(new_n1259), .C1(G107), .C2(new_n814), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n833), .A2(G97), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n818), .A2(new_n652), .B1(new_n1021), .B2(G77), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n820), .A2(G116), .B1(new_n804), .B2(G294), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n817), .A2(new_n202), .B1(new_n819), .B2(new_n1145), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n269), .B(new_n1265), .C1(G58), .C2(new_n1021), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n823), .A2(G137), .B1(new_n824), .B2(G128), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1266), .B(new_n1267), .C1(new_n1051), .C2(new_n813), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n804), .A2(G132), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT119), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n808), .B2(new_n834), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1264), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n876), .B(new_n1258), .C1(new_n1272), .C2(new_n794), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1257), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1252), .B2(new_n776), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1256), .A2(new_n1276), .ZN(G381));
  AOI21_X1  g1077(.A(new_n1249), .B1(new_n1210), .B2(new_n1218), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1183), .ZN(new_n1279));
  OR3_X1    g1079(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(G381), .A2(G387), .A3(G390), .A4(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1281), .B2(KEYINPUT120), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(KEYINPUT120), .B2(new_n1281), .ZN(G407));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(G343), .C2(new_n1279), .ZN(G409));
  INV_X1    g1084(.A(G390), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT125), .B1(G387), .B2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(new_n842), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1014), .B2(new_n1040), .ZN(new_n1289));
  AND3_X1   g1089(.A1(G390), .A2(new_n1014), .A3(new_n1040), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n1286), .A2(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G387), .A2(new_n1285), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G390), .A2(new_n1014), .A3(new_n1040), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1293), .A2(KEYINPUT125), .A3(new_n1294), .A4(new_n1287), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1291), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1183), .B1(new_n1219), .B2(new_n1250), .ZN(new_n1297));
  INV_X1    g1097(.A(G213), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1298), .A2(G343), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1175), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1254), .B(new_n1301), .C1(new_n1302), .C2(new_n1186), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1176), .A2(new_n1182), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1158), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT121), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n776), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(new_n1247), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1220), .A2(KEYINPUT121), .A3(new_n1248), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1300), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1253), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1252), .A2(KEYINPUT60), .A3(new_n1186), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n733), .A3(new_n1315), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT122), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n853), .B2(new_n879), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1316), .A2(new_n1276), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n734), .B1(new_n1313), .B2(new_n1253), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1275), .B1(new_n1323), .B2(new_n1315), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1324), .B2(new_n1319), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1297), .A2(new_n1312), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1296), .B1(new_n1326), .B2(KEYINPUT63), .ZN(new_n1327));
  XOR2_X1   g1127(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1328));
  NAND4_X1  g1128(.A1(new_n1183), .A2(new_n1303), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1329), .B(new_n1300), .C1(new_n1278), .C2(new_n1183), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1330), .B2(new_n1325), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1299), .A2(G2897), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1275), .B(new_n1320), .C1(new_n1323), .C2(new_n1315), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1319), .B1(new_n1316), .B2(new_n1276), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1332), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1322), .B(new_n1336), .C1(new_n1324), .C2(new_n1319), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1330), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(KEYINPUT124), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1330), .A2(new_n1338), .A3(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1327), .A2(new_n1331), .A3(new_n1340), .A4(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT61), .B1(new_n1330), .B2(new_n1338), .ZN(new_n1344));
  OAI21_X1  g1144(.A(KEYINPUT62), .B1(new_n1330), .B2(new_n1325), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1312), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(G375), .A2(G378), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT62), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1325), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1346), .A2(new_n1347), .A3(new_n1348), .A4(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1344), .A2(new_n1345), .A3(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT126), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1291), .A2(new_n1352), .A3(new_n1295), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1352), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1351), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1343), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1343), .A2(new_n1356), .A3(KEYINPUT127), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(G405));
  NAND2_X1  g1161(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1362), .B(new_n1325), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1347), .A2(new_n1279), .ZN(new_n1364));
  XNOR2_X1  g1164(.A(new_n1363), .B(new_n1364), .ZN(G402));
endmodule


