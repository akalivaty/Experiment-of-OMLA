

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732;

  OR2_X1 U372 ( .A1(n609), .A2(n421), .ZN(n426) );
  INV_X1 U373 ( .A(G953), .ZN(n705) );
  OR2_X1 U374 ( .A1(n511), .A2(n627), .ZN(n539) );
  OR2_X1 U375 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U376 ( .A(n372), .B(n371), .ZN(n647) );
  XNOR2_X1 U377 ( .A(n426), .B(n425), .ZN(n479) );
  OR2_X1 U378 ( .A1(n693), .A2(G902), .ZN(n389) );
  NOR2_X1 U379 ( .A1(n505), .A2(n571), .ZN(n507) );
  XNOR2_X1 U380 ( .A(n504), .B(KEYINPUT95), .ZN(n505) );
  INV_X1 U381 ( .A(KEYINPUT106), .ZN(n552) );
  NAND2_X1 U382 ( .A1(n668), .A2(n667), .ZN(n553) );
  XNOR2_X1 U383 ( .A(n487), .B(KEYINPUT0), .ZN(n498) );
  XNOR2_X1 U384 ( .A(n550), .B(n549), .ZN(n710) );
  XNOR2_X1 U385 ( .A(n529), .B(n528), .ZN(n682) );
  BUF_X1 U386 ( .A(n498), .Z(n501) );
  XNOR2_X1 U387 ( .A(n458), .B(n457), .ZN(n488) );
  XNOR2_X1 U388 ( .A(n606), .B(n605), .ZN(n704) );
  XOR2_X1 U389 ( .A(n581), .B(KEYINPUT80), .Z(n351) );
  XOR2_X1 U390 ( .A(n392), .B(KEYINPUT73), .Z(n352) );
  OR2_X1 U391 ( .A1(n589), .A2(KEYINPUT47), .ZN(n353) );
  OR2_X1 U392 ( .A1(n485), .A2(n484), .ZN(n354) );
  XOR2_X1 U393 ( .A(KEYINPUT3), .B(G119), .Z(n355) );
  NOR2_X1 U394 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U395 ( .A1(n540), .A2(n519), .ZN(n520) );
  INV_X1 U396 ( .A(KEYINPUT99), .ZN(n506) );
  XNOR2_X1 U397 ( .A(n398), .B(n397), .ZN(n399) );
  NOR2_X1 U398 ( .A1(n539), .A2(n538), .ZN(n548) );
  OR2_X1 U399 ( .A1(n647), .A2(n648), .ZN(n524) );
  XNOR2_X1 U400 ( .A(n400), .B(n399), .ZN(n618) );
  XNOR2_X1 U401 ( .A(n553), .B(n552), .ZN(n663) );
  XNOR2_X1 U402 ( .A(KEYINPUT98), .B(G478), .ZN(n457) );
  NOR2_X2 U403 ( .A1(n688), .A2(n599), .ZN(n690) );
  XNOR2_X1 U404 ( .A(n481), .B(n480), .ZN(n577) );
  BUF_X1 U405 ( .A(n690), .Z(n700) );
  XNOR2_X1 U406 ( .A(n555), .B(n554), .ZN(n681) );
  BUF_X1 U407 ( .A(n577), .Z(n587) );
  OR2_X1 U408 ( .A1(n489), .A2(n532), .ZN(n661) );
  XNOR2_X1 U409 ( .A(n497), .B(KEYINPUT32), .ZN(n518) );
  XNOR2_X1 U410 ( .A(n516), .B(KEYINPUT100), .ZN(n626) );
  INV_X1 U411 ( .A(KEYINPUT67), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n356), .B(KEYINPUT10), .ZN(n357) );
  XNOR2_X2 U413 ( .A(G146), .B(G125), .ZN(n416) );
  XNOR2_X2 U414 ( .A(n357), .B(n416), .ZN(n720) );
  XOR2_X1 U415 ( .A(KEYINPUT24), .B(G110), .Z(n359) );
  XNOR2_X1 U416 ( .A(G119), .B(G128), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n720), .B(n360), .ZN(n362) );
  XOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n368) );
  XNOR2_X1 U421 ( .A(G140), .B(G137), .ZN(n378) );
  XNOR2_X1 U422 ( .A(n378), .B(KEYINPUT74), .ZN(n366) );
  XOR2_X1 U423 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n364) );
  NAND2_X1 U424 ( .A1(G234), .A2(n705), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n454) );
  NAND2_X1 U426 ( .A1(G221), .A2(n454), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n701) );
  NOR2_X1 U429 ( .A1(n701), .A2(G902), .ZN(n372) );
  XNOR2_X1 U430 ( .A(KEYINPUT15), .B(G902), .ZN(n599) );
  NAND2_X1 U431 ( .A1(G234), .A2(n599), .ZN(n369) );
  XNOR2_X1 U432 ( .A(KEYINPUT20), .B(n369), .ZN(n373) );
  AND2_X1 U433 ( .A1(n373), .A2(G217), .ZN(n370) );
  XNOR2_X1 U434 ( .A(KEYINPUT25), .B(n370), .ZN(n371) );
  AND2_X1 U435 ( .A1(n373), .A2(G221), .ZN(n375) );
  INV_X1 U436 ( .A(KEYINPUT21), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n648) );
  INV_X1 U438 ( .A(n524), .ZN(n643) );
  XNOR2_X2 U439 ( .A(G143), .B(G128), .ZN(n449) );
  XNOR2_X1 U440 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n449), .B(n376), .ZN(n412) );
  INV_X1 U442 ( .A(G134), .ZN(n467) );
  XNOR2_X1 U443 ( .A(n467), .B(G131), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n412), .B(n377), .ZN(n398) );
  INV_X1 U445 ( .A(n398), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n379), .B(n378), .ZN(n719) );
  NAND2_X1 U447 ( .A1(n705), .A2(G227), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n380), .B(KEYINPUT75), .ZN(n381) );
  XNOR2_X1 U449 ( .A(KEYINPUT71), .B(G110), .ZN(n411) );
  XNOR2_X1 U450 ( .A(n381), .B(n411), .ZN(n385) );
  XNOR2_X1 U451 ( .A(G146), .B(G104), .ZN(n383) );
  XNOR2_X1 U452 ( .A(G101), .B(G107), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n719), .B(n386), .ZN(n693) );
  INV_X1 U456 ( .A(KEYINPUT69), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n387), .B(G469), .ZN(n388) );
  XNOR2_X2 U458 ( .A(n389), .B(n388), .ZN(n559) );
  NAND2_X1 U459 ( .A1(n643), .A2(n559), .ZN(n502) );
  XNOR2_X1 U460 ( .A(n502), .B(KEYINPUT104), .ZN(n405) );
  XOR2_X1 U461 ( .A(G116), .B(KEYINPUT5), .Z(n391) );
  NOR2_X1 U462 ( .A1(G953), .A2(G237), .ZN(n433) );
  NAND2_X1 U463 ( .A1(n433), .A2(G210), .ZN(n390) );
  XNOR2_X1 U464 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U465 ( .A(G137), .B(G146), .ZN(n393) );
  XNOR2_X1 U466 ( .A(n352), .B(n393), .ZN(n400) );
  XNOR2_X1 U467 ( .A(G113), .B(G101), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n355), .B(n394), .ZN(n396) );
  INV_X1 U469 ( .A(KEYINPUT70), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n408) );
  BUF_X1 U471 ( .A(n408), .Z(n397) );
  INV_X1 U472 ( .A(G902), .ZN(n437) );
  NAND2_X1 U473 ( .A1(n618), .A2(n437), .ZN(n401) );
  XNOR2_X2 U474 ( .A(n401), .B(G472), .ZN(n653) );
  INV_X1 U475 ( .A(G237), .ZN(n402) );
  NAND2_X1 U476 ( .A1(n437), .A2(n402), .ZN(n422) );
  NAND2_X1 U477 ( .A1(n422), .A2(G214), .ZN(n667) );
  NAND2_X1 U478 ( .A1(n653), .A2(n667), .ZN(n403) );
  XNOR2_X1 U479 ( .A(n403), .B(KEYINPUT30), .ZN(n404) );
  NOR2_X1 U480 ( .A1(n405), .A2(n404), .ZN(n464) );
  XOR2_X2 U481 ( .A(G116), .B(G107), .Z(n448) );
  XOR2_X1 U482 ( .A(KEYINPUT72), .B(KEYINPUT16), .Z(n406) );
  XNOR2_X1 U483 ( .A(n448), .B(n406), .ZN(n407) );
  XOR2_X1 U484 ( .A(G122), .B(G104), .Z(n427) );
  XNOR2_X1 U485 ( .A(n407), .B(n427), .ZN(n409) );
  XNOR2_X1 U486 ( .A(n409), .B(n408), .ZN(n706) );
  XNOR2_X1 U487 ( .A(KEYINPUT76), .B(KEYINPUT89), .ZN(n410) );
  XNOR2_X1 U488 ( .A(n411), .B(n410), .ZN(n413) );
  XNOR2_X1 U489 ( .A(n413), .B(n412), .ZN(n419) );
  XNOR2_X1 U490 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n415) );
  NAND2_X1 U491 ( .A1(n705), .A2(G224), .ZN(n414) );
  XNOR2_X1 U492 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U493 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U494 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U495 ( .A(n706), .B(n420), .ZN(n609) );
  INV_X1 U496 ( .A(n599), .ZN(n421) );
  NAND2_X1 U497 ( .A1(n422), .A2(G210), .ZN(n424) );
  INV_X1 U498 ( .A(KEYINPUT90), .ZN(n423) );
  XNOR2_X1 U499 ( .A(n424), .B(n423), .ZN(n425) );
  BUF_X1 U500 ( .A(n479), .Z(n462) );
  INV_X1 U501 ( .A(n462), .ZN(n565) );
  XNOR2_X1 U502 ( .A(G113), .B(G143), .ZN(n428) );
  XNOR2_X1 U503 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U504 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n430) );
  XNOR2_X1 U505 ( .A(G131), .B(G140), .ZN(n429) );
  XNOR2_X1 U506 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U507 ( .A(n432), .B(n431), .Z(n436) );
  AND2_X1 U508 ( .A1(G214), .A2(n433), .ZN(n434) );
  XNOR2_X1 U509 ( .A(n720), .B(n434), .ZN(n435) );
  XNOR2_X1 U510 ( .A(n436), .B(n435), .ZN(n601) );
  NAND2_X1 U511 ( .A1(n601), .A2(n437), .ZN(n439) );
  XNOR2_X1 U512 ( .A(KEYINPUT13), .B(G475), .ZN(n438) );
  XNOR2_X1 U513 ( .A(n439), .B(n438), .ZN(n489) );
  INV_X1 U514 ( .A(n489), .ZN(n533) );
  NAND2_X1 U515 ( .A1(G234), .A2(G237), .ZN(n440) );
  XNOR2_X1 U516 ( .A(n440), .B(KEYINPUT14), .ZN(n444) );
  NAND2_X1 U517 ( .A1(G902), .A2(n444), .ZN(n441) );
  XNOR2_X1 U518 ( .A(KEYINPUT91), .B(n441), .ZN(n442) );
  NAND2_X1 U519 ( .A1(n442), .A2(G953), .ZN(n482) );
  XNOR2_X1 U520 ( .A(KEYINPUT102), .B(n482), .ZN(n443) );
  NOR2_X1 U521 ( .A1(G900), .A2(n443), .ZN(n445) );
  NAND2_X1 U522 ( .A1(G952), .A2(n444), .ZN(n680) );
  NOR2_X1 U523 ( .A1(n680), .A2(G953), .ZN(n484) );
  NOR2_X1 U524 ( .A1(n445), .A2(n484), .ZN(n471) );
  XOR2_X1 U525 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n447) );
  XNOR2_X1 U526 ( .A(G134), .B(G122), .ZN(n446) );
  XNOR2_X1 U527 ( .A(n447), .B(n446), .ZN(n453) );
  XNOR2_X1 U528 ( .A(KEYINPUT96), .B(KEYINPUT9), .ZN(n450) );
  XNOR2_X1 U529 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U530 ( .A(n448), .B(n451), .ZN(n452) );
  XOR2_X1 U531 ( .A(n453), .B(n452), .Z(n456) );
  NAND2_X1 U532 ( .A1(G217), .A2(n454), .ZN(n455) );
  XNOR2_X1 U533 ( .A(n456), .B(n455), .ZN(n697) );
  NOR2_X1 U534 ( .A1(G902), .A2(n697), .ZN(n458) );
  NOR2_X1 U535 ( .A1(n471), .A2(n488), .ZN(n459) );
  NAND2_X1 U536 ( .A1(n533), .A2(n459), .ZN(n460) );
  NOR2_X1 U537 ( .A1(n565), .A2(n460), .ZN(n461) );
  NAND2_X1 U538 ( .A1(n464), .A2(n461), .ZN(n573) );
  XNOR2_X1 U539 ( .A(n573), .B(G143), .ZN(G45) );
  XNOR2_X1 U540 ( .A(n462), .B(KEYINPUT38), .ZN(n551) );
  NOR2_X1 U541 ( .A1(n551), .A2(n471), .ZN(n463) );
  NAND2_X1 U542 ( .A1(n464), .A2(n463), .ZN(n466) );
  XNOR2_X1 U543 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n465) );
  XNOR2_X1 U544 ( .A(n466), .B(n465), .ZN(n468) );
  INV_X1 U545 ( .A(n488), .ZN(n532) );
  NAND2_X1 U546 ( .A1(n489), .A2(n532), .ZN(n662) );
  NOR2_X1 U547 ( .A1(n468), .A2(n662), .ZN(n594) );
  XNOR2_X1 U548 ( .A(n594), .B(n467), .ZN(G36) );
  NOR2_X1 U549 ( .A1(n468), .A2(n661), .ZN(n470) );
  XOR2_X1 U550 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n469) );
  XNOR2_X1 U551 ( .A(n470), .B(n469), .ZN(n562) );
  XOR2_X1 U552 ( .A(G131), .B(n562), .Z(G33) );
  NOR2_X1 U553 ( .A1(n648), .A2(n471), .ZN(n472) );
  XNOR2_X1 U554 ( .A(KEYINPUT68), .B(n472), .ZN(n473) );
  NAND2_X1 U555 ( .A1(n473), .A2(n647), .ZN(n556) );
  XNOR2_X1 U556 ( .A(n653), .B(KEYINPUT6), .ZN(n525) );
  NOR2_X1 U557 ( .A1(n556), .A2(n525), .ZN(n474) );
  XNOR2_X1 U558 ( .A(n474), .B(KEYINPUT103), .ZN(n475) );
  NOR2_X1 U559 ( .A1(n661), .A2(n475), .ZN(n476) );
  NAND2_X1 U560 ( .A1(n476), .A2(n667), .ZN(n566) );
  XNOR2_X2 U561 ( .A(n559), .B(KEYINPUT1), .ZN(n642) );
  NOR2_X1 U562 ( .A1(n566), .A2(n642), .ZN(n477) );
  XNOR2_X1 U563 ( .A(n477), .B(KEYINPUT43), .ZN(n478) );
  NOR2_X1 U564 ( .A1(n478), .A2(n462), .ZN(n595) );
  XOR2_X1 U565 ( .A(G140), .B(n595), .Z(G42) );
  NAND2_X1 U566 ( .A1(n479), .A2(n667), .ZN(n481) );
  INV_X1 U567 ( .A(KEYINPUT19), .ZN(n480) );
  INV_X1 U568 ( .A(n577), .ZN(n486) );
  NOR2_X1 U569 ( .A1(G898), .A2(n482), .ZN(n483) );
  XNOR2_X1 U570 ( .A(n483), .B(KEYINPUT92), .ZN(n485) );
  NAND2_X1 U571 ( .A1(n486), .A2(n354), .ZN(n487) );
  AND2_X1 U572 ( .A1(n489), .A2(n488), .ZN(n666) );
  INV_X1 U573 ( .A(n648), .ZN(n490) );
  NAND2_X1 U574 ( .A1(n666), .A2(n490), .ZN(n491) );
  OR2_X2 U575 ( .A1(n498), .A2(n491), .ZN(n493) );
  INV_X1 U576 ( .A(KEYINPUT22), .ZN(n492) );
  XNOR2_X2 U577 ( .A(n493), .B(n492), .ZN(n515) );
  AND2_X1 U578 ( .A1(n525), .A2(n647), .ZN(n494) );
  NAND2_X1 U579 ( .A1(n494), .A2(n642), .ZN(n495) );
  XNOR2_X1 U580 ( .A(n495), .B(KEYINPUT77), .ZN(n496) );
  NAND2_X1 U581 ( .A1(n515), .A2(n496), .ZN(n497) );
  XNOR2_X1 U582 ( .A(n518), .B(G119), .ZN(G21) );
  INV_X1 U583 ( .A(n653), .ZN(n557) );
  NOR2_X1 U584 ( .A1(n524), .A2(n557), .ZN(n499) );
  NAND2_X1 U585 ( .A1(n499), .A2(n642), .ZN(n656) );
  NOR2_X1 U586 ( .A1(n501), .A2(n656), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n500), .B(KEYINPUT31), .ZN(n640) );
  XNOR2_X1 U588 ( .A(n501), .B(KEYINPUT93), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n502), .A2(n653), .ZN(n503) );
  NAND2_X1 U590 ( .A1(n530), .A2(n503), .ZN(n629) );
  NAND2_X1 U591 ( .A1(n640), .A2(n629), .ZN(n504) );
  AND2_X1 U592 ( .A1(n662), .A2(n661), .ZN(n571) );
  XNOR2_X1 U593 ( .A(n507), .B(n506), .ZN(n511) );
  INV_X1 U594 ( .A(n647), .ZN(n508) );
  NAND2_X1 U595 ( .A1(n525), .A2(n508), .ZN(n509) );
  NOR2_X1 U596 ( .A1(n509), .A2(n642), .ZN(n510) );
  AND2_X1 U597 ( .A1(n515), .A2(n510), .ZN(n627) );
  AND2_X1 U598 ( .A1(n557), .A2(n647), .ZN(n513) );
  INV_X1 U599 ( .A(n642), .ZN(n512) );
  AND2_X1 U600 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U601 ( .A1(n515), .A2(n514), .ZN(n516) );
  AND2_X1 U602 ( .A1(n626), .A2(n518), .ZN(n517) );
  NOR2_X1 U603 ( .A1(n517), .A2(KEYINPUT85), .ZN(n521) );
  NAND2_X1 U604 ( .A1(n518), .A2(n626), .ZN(n540) );
  NOR2_X1 U605 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n519) );
  NOR2_X1 U606 ( .A1(n521), .A2(n520), .ZN(n523) );
  INV_X1 U607 ( .A(KEYINPUT84), .ZN(n522) );
  NOR2_X1 U608 ( .A1(n523), .A2(n522), .ZN(n537) );
  NOR2_X1 U609 ( .A1(n525), .A2(n524), .ZN(n526) );
  AND2_X1 U610 ( .A1(n526), .A2(n642), .ZN(n529) );
  XNOR2_X1 U611 ( .A(KEYINPUT101), .B(KEYINPUT33), .ZN(n527) );
  XNOR2_X1 U612 ( .A(n527), .B(KEYINPUT86), .ZN(n528) );
  NAND2_X1 U613 ( .A1(n530), .A2(n682), .ZN(n531) );
  XNOR2_X1 U614 ( .A(n531), .B(KEYINPUT34), .ZN(n535) );
  NAND2_X1 U615 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U616 ( .A(n536), .B(KEYINPUT35), .ZN(n625) );
  NOR2_X1 U617 ( .A1(n537), .A2(n625), .ZN(n538) );
  NAND2_X1 U618 ( .A1(n625), .A2(KEYINPUT84), .ZN(n543) );
  INV_X1 U619 ( .A(n540), .ZN(n541) );
  AND2_X1 U620 ( .A1(n541), .A2(KEYINPUT44), .ZN(n542) );
  NAND2_X1 U621 ( .A1(n543), .A2(n542), .ZN(n546) );
  INV_X1 U622 ( .A(KEYINPUT44), .ZN(n544) );
  NAND2_X1 U623 ( .A1(n544), .A2(KEYINPUT84), .ZN(n545) );
  NAND2_X1 U624 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U625 ( .A1(n548), .A2(n547), .ZN(n550) );
  XOR2_X1 U626 ( .A(KEYINPUT82), .B(KEYINPUT45), .Z(n549) );
  INV_X1 U627 ( .A(n551), .ZN(n668) );
  NAND2_X1 U628 ( .A1(n666), .A2(n663), .ZN(n555) );
  XNOR2_X1 U629 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n554) );
  NOR2_X1 U630 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U631 ( .A(KEYINPUT28), .B(n558), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n560), .A2(n559), .ZN(n582) );
  NOR2_X1 U633 ( .A1(n681), .A2(n582), .ZN(n561) );
  XNOR2_X1 U634 ( .A(n561), .B(KEYINPUT42), .ZN(n732) );
  NOR2_X1 U635 ( .A1(n732), .A2(n562), .ZN(n564) );
  XNOR2_X1 U636 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n563) );
  XNOR2_X1 U637 ( .A(n564), .B(n563), .ZN(n592) );
  XOR2_X1 U638 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n568) );
  NOR2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U640 ( .A(n568), .B(n567), .Z(n569) );
  NAND2_X1 U641 ( .A1(n569), .A2(n642), .ZN(n570) );
  XNOR2_X1 U642 ( .A(n570), .B(KEYINPUT109), .ZN(n730) );
  NAND2_X1 U643 ( .A1(KEYINPUT47), .A2(n571), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT81), .ZN(n575) );
  INV_X1 U645 ( .A(n573), .ZN(n574) );
  XNOR2_X1 U646 ( .A(KEYINPUT78), .B(n576), .ZN(n580) );
  OR2_X1 U647 ( .A1(n582), .A2(n587), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n578), .A2(KEYINPUT47), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U650 ( .A(n582), .ZN(n586) );
  INV_X1 U651 ( .A(n662), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n586), .A2(n583), .ZN(n584) );
  NOR2_X1 U653 ( .A1(n584), .A2(n587), .ZN(n633) );
  INV_X1 U654 ( .A(n661), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n588) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n636) );
  NOR2_X1 U657 ( .A1(n633), .A2(n636), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n351), .A2(n353), .ZN(n590) );
  NOR2_X1 U659 ( .A1(n730), .A2(n590), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U661 ( .A(KEYINPUT48), .B(n593), .Z(n597) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n721) );
  NOR2_X1 U664 ( .A1(n710), .A2(n721), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT2), .ZN(n688) );
  NAND2_X1 U666 ( .A1(n690), .A2(G475), .ZN(n603) );
  XOR2_X1 U667 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n600) );
  XNOR2_X1 U668 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n603), .B(n602), .ZN(n607) );
  INV_X1 U670 ( .A(G952), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n604), .A2(G953), .ZN(n606) );
  INV_X1 U672 ( .A(KEYINPUT88), .ZN(n605) );
  NOR2_X1 U673 ( .A1(n607), .A2(n704), .ZN(n608) );
  XNOR2_X1 U674 ( .A(n608), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U675 ( .A1(n690), .A2(G210), .ZN(n614) );
  BUF_X1 U676 ( .A(n609), .Z(n612) );
  XNOR2_X1 U677 ( .A(KEYINPUT79), .B(KEYINPUT54), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n610), .B(KEYINPUT55), .ZN(n611) );
  XNOR2_X1 U679 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U680 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X1 U681 ( .A1(n615), .A2(n704), .ZN(n617) );
  XOR2_X1 U682 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n616) );
  XNOR2_X1 U683 ( .A(n617), .B(n616), .ZN(G51) );
  NAND2_X1 U684 ( .A1(n690), .A2(G472), .ZN(n621) );
  XOR2_X1 U685 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n619) );
  XNOR2_X1 U686 ( .A(n618), .B(n619), .ZN(n620) );
  XNOR2_X1 U687 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n622), .A2(n704), .ZN(n624) );
  XNOR2_X1 U689 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n623) );
  XNOR2_X1 U690 ( .A(n624), .B(n623), .ZN(G57) );
  XOR2_X1 U691 ( .A(G122), .B(n625), .Z(G24) );
  XNOR2_X1 U692 ( .A(n626), .B(G110), .ZN(G12) );
  XOR2_X1 U693 ( .A(G101), .B(n627), .Z(G3) );
  NOR2_X1 U694 ( .A1(n661), .A2(n629), .ZN(n628) );
  XOR2_X1 U695 ( .A(G104), .B(n628), .Z(G6) );
  NOR2_X1 U696 ( .A1(n662), .A2(n629), .ZN(n631) );
  XNOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U699 ( .A(G107), .B(n632), .ZN(G9) );
  XOR2_X1 U700 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n635) );
  XNOR2_X1 U701 ( .A(G128), .B(n633), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n635), .B(n634), .ZN(G30) );
  XOR2_X1 U703 ( .A(G146), .B(n636), .Z(n637) );
  XNOR2_X1 U704 ( .A(KEYINPUT112), .B(n637), .ZN(G48) );
  NOR2_X1 U705 ( .A1(n661), .A2(n640), .ZN(n639) );
  XNOR2_X1 U706 ( .A(G113), .B(KEYINPUT113), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(G15) );
  NOR2_X1 U708 ( .A1(n662), .A2(n640), .ZN(n641) );
  XOR2_X1 U709 ( .A(G116), .B(n641), .Z(G18) );
  NOR2_X1 U710 ( .A1(n643), .A2(n642), .ZN(n645) );
  XNOR2_X1 U711 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n646), .B(KEYINPUT116), .ZN(n655) );
  XOR2_X1 U714 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n650) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT114), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U720 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U721 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NOR2_X1 U722 ( .A1(n681), .A2(n659), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT118), .ZN(n676) );
  NAND2_X1 U724 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U726 ( .A(n665), .B(KEYINPUT119), .ZN(n672) );
  INV_X1 U727 ( .A(n666), .ZN(n670) );
  NOR2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n674) );
  INV_X1 U731 ( .A(n682), .ZN(n673) );
  NOR2_X1 U732 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U733 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  XNOR2_X1 U735 ( .A(KEYINPUT120), .B(n678), .ZN(n679) );
  NOR2_X1 U736 ( .A1(n680), .A2(n679), .ZN(n686) );
  INV_X1 U737 ( .A(n681), .ZN(n683) );
  NAND2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U739 ( .A1(n684), .A2(n705), .ZN(n685) );
  NOR2_X1 U740 ( .A1(n686), .A2(n685), .ZN(n687) );
  AND2_X1 U741 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n689), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U743 ( .A1(n700), .A2(G469), .ZN(n695) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U745 ( .A(n691), .B(KEYINPUT122), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U747 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U748 ( .A1(n704), .A2(n696), .ZN(G54) );
  NAND2_X1 U749 ( .A1(n700), .A2(G478), .ZN(n698) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U751 ( .A1(n704), .A2(n699), .ZN(G63) );
  NAND2_X1 U752 ( .A1(n700), .A2(G217), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U754 ( .A1(n704), .A2(n703), .ZN(G66) );
  NOR2_X1 U755 ( .A1(G898), .A2(n705), .ZN(n709) );
  BUF_X1 U756 ( .A(n706), .Z(n707) );
  XOR2_X1 U757 ( .A(n707), .B(G110), .Z(n708) );
  NOR2_X1 U758 ( .A1(n709), .A2(n708), .ZN(n718) );
  NOR2_X1 U759 ( .A1(n710), .A2(G953), .ZN(n711) );
  XNOR2_X1 U760 ( .A(n711), .B(KEYINPUT125), .ZN(n716) );
  NAND2_X1 U761 ( .A1(G224), .A2(G953), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n712), .B(KEYINPUT61), .ZN(n713) );
  XNOR2_X1 U763 ( .A(KEYINPUT124), .B(n713), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U767 ( .A(n720), .B(n719), .Z(n723) );
  XNOR2_X1 U768 ( .A(n721), .B(n723), .ZN(n722) );
  NOR2_X1 U769 ( .A1(n722), .A2(G953), .ZN(n728) );
  XOR2_X1 U770 ( .A(G227), .B(n723), .Z(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n725), .A2(G953), .ZN(n726) );
  XOR2_X1 U773 ( .A(KEYINPUT126), .B(n726), .Z(n727) );
  NOR2_X1 U774 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U775 ( .A(KEYINPUT127), .B(n729), .ZN(G72) );
  XNOR2_X1 U776 ( .A(G125), .B(n730), .ZN(n731) );
  XNOR2_X1 U777 ( .A(n731), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U778 ( .A(G137), .B(n732), .Z(G39) );
endmodule

