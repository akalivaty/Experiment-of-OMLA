//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208));
  NOR4_X1   g007(.A1(new_n208), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT89), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n207), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT90), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G43gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G50gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT88), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G29gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n211), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT15), .B1(new_n216), .B2(new_n218), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n219), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(new_n207), .C1(new_n209), .C2(new_n212), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n214), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n211), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n219), .B(new_n230), .C1(new_n224), .C2(new_n207), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G15gat), .B(G22gat), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT16), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(G1gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G8gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n238), .A2(new_n239), .A3(G8gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT17), .A3(new_n231), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n234), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n232), .B1(new_n242), .B2(new_n243), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n248), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n247), .B(KEYINPUT13), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n244), .A2(new_n231), .A3(new_n229), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n248), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AND4_X1   g056(.A1(new_n206), .A2(new_n251), .A3(new_n252), .A4(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n249), .B2(new_n250), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n206), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(new_n252), .A3(new_n257), .ZN(new_n263));
  INV_X1    g062(.A(new_n206), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n259), .A2(new_n206), .A3(new_n252), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT91), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n269));
  XOR2_X1   g068(.A(G127gat), .B(G134gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(KEYINPUT1), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT67), .ZN(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT1), .B1(new_n271), .B2(KEYINPUT68), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(new_n277), .C1(KEYINPUT68), .C2(new_n271), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT2), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G148gat), .ZN(new_n283));
  INV_X1    g082(.A(G148gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G141gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n281), .A2(KEYINPUT72), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(KEYINPUT72), .B2(new_n281), .ZN(new_n287));
  XOR2_X1   g086(.A(G155gat), .B(G162gat), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT73), .B(G148gat), .Z(new_n290));
  OAI21_X1  g089(.A(new_n283), .B1(new_n290), .B2(new_n282), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n291), .A2(new_n281), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n269), .B1(new_n279), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n281), .A3(new_n295), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n299), .A2(new_n291), .B1(new_n288), .B2(new_n287), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n300), .A2(KEYINPUT4), .A3(new_n273), .A4(new_n278), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n296), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(KEYINPUT3), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n307));
  AOI22_X1  g106(.A1(new_n300), .A2(new_n307), .B1(new_n273), .B2(new_n278), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT77), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n302), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT5), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n302), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n306), .A2(new_n311), .A3(new_n308), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n311), .B1(new_n306), .B2(new_n308), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n314), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n279), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n300), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n279), .A3(new_n305), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT5), .B1(new_n323), .B2(new_n314), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n315), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT85), .ZN(new_n327));
  XOR2_X1   g126(.A(G57gat), .B(G85gat), .Z(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT79), .ZN(new_n329));
  XOR2_X1   g128(.A(G1gat), .B(G29gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n325), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT6), .B1(new_n326), .B2(new_n333), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n315), .A2(new_n325), .A3(KEYINPUT6), .A4(new_n334), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT22), .ZN(new_n345));
  INV_X1    g144(.A(G211gat), .ZN(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT71), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  INV_X1    g152(.A(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G183gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n354), .ZN(new_n359));
  NOR2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n360), .A2(KEYINPUT26), .ZN(new_n361));
  INV_X1    g160(.A(new_n360), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  AOI211_X1 g162(.A(new_n359), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n365));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n359), .A2(KEYINPUT24), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n358), .A2(new_n354), .ZN(new_n373));
  NAND3_X1  g172(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n374), .A2(KEYINPUT64), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(KEYINPUT64), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n357), .A2(new_n364), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n373), .B(KEYINPUT66), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n374), .B1(new_n380), .B2(new_n359), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n369), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT25), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  INV_X1    g183(.A(G226gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n378), .A2(new_n383), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n378), .A2(new_n383), .A3(new_n388), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n352), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n391), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n349), .B(new_n350), .Z(new_n394));
  NOR3_X1   g193(.A1(new_n393), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n343), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT37), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n390), .B2(new_n391), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399));
  INV_X1    g198(.A(new_n352), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(new_n391), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n399), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n392), .B2(new_n395), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT38), .ZN(new_n406));
  INV_X1    g205(.A(new_n343), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n396), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n351), .A3(new_n391), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n400), .B1(new_n393), .B2(new_n389), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT37), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n407), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(KEYINPUT87), .A3(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n405), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n409), .B1(new_n417), .B2(KEYINPUT38), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n339), .A2(new_n340), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(new_n215), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n289), .A2(new_n296), .A3(new_n307), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n384), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n352), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n351), .A2(KEYINPUT29), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n303), .B(new_n305), .C1(KEYINPUT3), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n394), .A2(new_n384), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n300), .B1(new_n433), .B2(new_n307), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n394), .B1(new_n427), .B2(new_n384), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n424), .B1(new_n437), .B2(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n432), .A2(new_n442), .A3(new_n436), .A4(new_n439), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n438), .A2(new_n441), .A3(new_n446), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n437), .A2(G22gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n440), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n424), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n410), .A2(new_n411), .A3(new_n407), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n455), .B(new_n343), .C1(new_n392), .C2(new_n395), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n323), .B2(new_n314), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n313), .B2(new_n314), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n462));
  INV_X1    g261(.A(new_n314), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n461), .A2(KEYINPUT40), .A3(new_n333), .A4(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(new_n333), .A3(new_n465), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(KEYINPUT84), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT84), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n467), .B(new_n337), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n419), .A2(new_n452), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n378), .A2(new_n383), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n320), .ZN(new_n477));
  INV_X1    g276(.A(G227gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n386), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n279), .A2(new_n383), .A3(new_n378), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT32), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(G15gat), .B(G43gat), .Z(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n481), .B(KEYINPUT32), .C1(new_n483), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n477), .A2(new_n480), .ZN(new_n492));
  INV_X1    g291(.A(new_n479), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT34), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n491), .B1(new_n498), .B2(KEYINPUT70), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n497), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n500), .A2(new_n490), .A3(new_n488), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n475), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n491), .A2(new_n498), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n490), .A3(new_n488), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n503), .B1(new_n475), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n321), .A2(new_n322), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n463), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n313), .B2(new_n314), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n319), .A2(new_n508), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n333), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n315), .A2(new_n325), .A3(new_n334), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n340), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n457), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n445), .A2(new_n447), .B1(new_n450), .B2(new_n424), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n507), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n474), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT35), .B1(new_n339), .B2(new_n340), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n519), .A2(new_n506), .A3(new_n458), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n499), .A2(new_n502), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n517), .A2(new_n452), .A3(new_n457), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n268), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G190gat), .B(G218gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT94), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT95), .B1(new_n532), .B2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n536), .A2(new_n537), .A3(G85gat), .A4(G92gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n532), .A2(new_n539), .A3(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G99gat), .B(G106gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n541), .A2(new_n547), .A3(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n234), .A2(new_n245), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n541), .A2(new_n547), .A3(new_n545), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n547), .B1(new_n541), .B2(new_n545), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n232), .A2(new_n555), .B1(KEYINPUT41), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n531), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(KEYINPUT98), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  NOR2_X1   g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n552), .A2(new_n531), .A3(new_n557), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT96), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n552), .A2(new_n566), .A3(new_n531), .A4(new_n557), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n558), .A2(KEYINPUT98), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n565), .A2(new_n571), .A3(new_n567), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n565), .B2(new_n567), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n572), .A2(new_n573), .A3(new_n558), .ZN(new_n574));
  INV_X1    g373(.A(new_n562), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(G57gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT92), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G57gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n581), .A3(G64gat), .ZN(new_n582));
  INV_X1    g381(.A(G64gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(G57gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n578), .A2(G64gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT9), .ZN(new_n592));
  INV_X1    g391(.A(new_n586), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n593), .A2(new_n588), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n585), .A2(new_n589), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n244), .B1(new_n597), .B2(new_n596), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n605), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n577), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n547), .A2(KEYINPUT99), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n549), .A2(new_n550), .A3(new_n595), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n592), .A2(new_n594), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n582), .A2(new_n584), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n587), .A2(new_n588), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n619), .B(new_n617), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n553), .B2(new_n554), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n555), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n616), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n615), .B1(new_n618), .B2(new_n623), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n614), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n626), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n630), .B2(new_n615), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT100), .B1(new_n631), .B2(new_n613), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633));
  NOR4_X1   g432(.A1(new_n627), .A2(new_n633), .A3(new_n628), .A4(new_n614), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n629), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n629), .B(KEYINPUT101), .C1(new_n632), .C2(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n610), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n529), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n517), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n236), .ZN(G1324gat));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n241), .B1(new_n644), .B2(new_n458), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT16), .B(G8gat), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n641), .A2(new_n457), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(KEYINPUT42), .B2(new_n647), .ZN(G1325gat));
  NAND2_X1  g448(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n504), .A2(new_n475), .A3(new_n505), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(G15gat), .B1(new_n641), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n506), .A2(G15gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n641), .B2(new_n654), .ZN(G1326gat));
  NOR2_X1   g454(.A1(new_n641), .A2(new_n452), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT43), .B(G22gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  NAND2_X1  g457(.A1(new_n221), .A2(new_n223), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n577), .B1(new_n521), .B2(new_n528), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT44), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(KEYINPUT44), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n609), .ZN(new_n664));
  INV_X1    g463(.A(new_n639), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n265), .A2(new_n266), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n659), .B1(new_n670), .B2(new_n517), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n666), .A2(new_n577), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n529), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(new_n517), .A3(new_n659), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(G1328gat));
  OAI21_X1  g476(.A(G36gat), .B1(new_n670), .B2(new_n457), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  AOI21_X1  g478(.A(G36gat), .B1(new_n679), .B2(KEYINPUT46), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n529), .A2(new_n458), .A3(new_n672), .A4(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(KEYINPUT46), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(new_n683), .ZN(G1329gat));
  OAI21_X1  g483(.A(new_n217), .B1(new_n673), .B2(new_n506), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n652), .A2(new_n217), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n670), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT47), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n690), .B(new_n685), .C1(new_n670), .C2(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(G1330gat));
  NOR3_X1   g491(.A1(new_n673), .A2(G50gat), .A3(new_n452), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n661), .A2(new_n519), .A3(new_n662), .A4(new_n669), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G50gat), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n694), .B2(G50gat), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI221_X4 g498(.A(new_n693), .B1(new_n696), .B2(KEYINPUT48), .C1(new_n694), .C2(G50gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(G1331gat));
  NAND2_X1  g500(.A1(new_n521), .A2(new_n528), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n610), .A2(new_n667), .A3(new_n665), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n517), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n579), .A2(new_n581), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1332gat));
  AOI21_X1  g507(.A(new_n457), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT105), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1333gat));
  INV_X1    g512(.A(new_n704), .ZN(new_n714));
  OAI21_X1  g513(.A(G71gat), .B1(new_n714), .B2(new_n652), .ZN(new_n715));
  INV_X1    g514(.A(G71gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n506), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n704), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n519), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT106), .B(G78gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n665), .A2(new_n609), .A3(new_n667), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n663), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n517), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n609), .A2(new_n667), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n458), .B1(new_n516), .B2(new_n340), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n652), .B1(new_n728), .B2(new_n452), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n458), .A2(new_n466), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n333), .B1(new_n326), .B2(KEYINPUT85), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n336), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n468), .A2(new_n469), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT84), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n470), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n519), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n729), .B1(new_n737), .B2(new_n419), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n523), .A2(new_n522), .B1(new_n526), .B2(KEYINPUT35), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n576), .B(new_n727), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n702), .A2(KEYINPUT51), .A3(new_n576), .A4(new_n727), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n705), .A2(new_n543), .A3(new_n639), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n726), .B1(new_n745), .B2(new_n746), .ZN(G1336gat));
  NAND3_X1  g546(.A1(new_n742), .A2(KEYINPUT108), .A3(new_n743), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n740), .A2(new_n749), .A3(new_n741), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n665), .A2(G92gat), .A3(new_n457), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT107), .Z(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n748), .A2(new_n750), .A3(new_n755), .A4(new_n752), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n661), .A2(new_n458), .A3(new_n662), .A4(new_n724), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G92gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n744), .A2(KEYINPUT110), .A3(new_n751), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT110), .B1(new_n744), .B2(new_n751), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n758), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1337gat));
  XNOR2_X1  g564(.A(KEYINPUT111), .B(G99gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n725), .B2(new_n652), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n717), .A2(new_n639), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n768), .A2(new_n766), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n745), .B2(new_n769), .ZN(G1338gat));
  NAND4_X1  g569(.A1(new_n661), .A2(new_n519), .A3(new_n662), .A4(new_n724), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n452), .A2(G106gat), .A3(new_n665), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n748), .A2(new_n750), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n744), .A2(new_n773), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n772), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1339gat));
  NAND2_X1  g579(.A1(new_n630), .A2(new_n615), .ZN(new_n781));
  INV_X1    g580(.A(new_n628), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(new_n613), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n633), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n631), .A2(KEYINPUT100), .A3(new_n613), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n613), .B1(new_n627), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(KEYINPUT54), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n625), .A2(new_n626), .A3(new_n616), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT55), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n790), .A2(new_n627), .A3(new_n787), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n630), .A2(new_n787), .A3(new_n615), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n614), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n786), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n667), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n248), .A2(new_n255), .A3(new_n254), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n205), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n266), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n637), .B2(new_n638), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n577), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n802), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n576), .A2(new_n805), .A3(new_n797), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n609), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n610), .A2(new_n667), .A3(new_n639), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n517), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n523), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT113), .Z(new_n812));
  INV_X1    g611(.A(G113gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(new_n268), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n452), .A2(new_n457), .A3(new_n525), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n667), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n814), .A2(new_n818), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n812), .B2(new_n665), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n665), .A2(G120gat), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT114), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n816), .B2(new_n822), .ZN(G1341gat));
  OAI21_X1  g622(.A(G127gat), .B1(new_n812), .B2(new_n664), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n664), .A2(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n816), .B2(new_n825), .ZN(G1342gat));
  OAI21_X1  g625(.A(G134gat), .B1(new_n812), .B2(new_n577), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n816), .A2(G134gat), .A3(new_n577), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT56), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1343gat));
  NOR3_X1   g629(.A1(new_n507), .A2(new_n517), .A3(new_n458), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  XOR2_X1   g631(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n793), .B2(new_n795), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n786), .A2(new_n791), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n262), .B2(new_n267), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n639), .A2(new_n805), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n261), .B1(new_n258), .B2(new_n260), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n265), .A2(KEYINPUT91), .A3(new_n266), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n803), .A3(KEYINPUT116), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n577), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n806), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n808), .B1(new_n845), .B2(new_n664), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n519), .A2(KEYINPUT57), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n809), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n849), .B2(new_n519), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n831), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n268), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n652), .A2(new_n519), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n457), .B1(new_n853), .B2(KEYINPUT117), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(KEYINPUT117), .B2(new_n853), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n810), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(G141gat), .A3(new_n268), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n851), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n667), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n857), .B1(new_n861), .B2(G141gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G1344gat));
  NOR3_X1   g663(.A1(new_n856), .A2(new_n290), .A3(new_n665), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n290), .B1(new_n851), .B2(new_n665), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n809), .A2(new_n847), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n558), .B1(new_n568), .B2(KEYINPUT97), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n565), .A2(new_n571), .A3(new_n567), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n575), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n570), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n870), .B(new_n797), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n805), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n870), .B1(new_n576), .B2(new_n797), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n844), .A2(new_n878), .A3(KEYINPUT119), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n837), .A2(new_n838), .A3(new_n832), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT116), .B1(new_n842), .B2(new_n803), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n576), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n876), .A2(new_n877), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n879), .A2(new_n885), .A3(new_n664), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n640), .A2(new_n268), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n452), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n869), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(new_n639), .A3(new_n831), .ZN(new_n890));
  NAND2_X1  g689(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n868), .B1(new_n890), .B2(new_n891), .ZN(G1345gat));
  INV_X1    g691(.A(new_n856), .ZN(new_n893));
  AOI21_X1  g692(.A(G155gat), .B1(new_n893), .B2(new_n609), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n609), .A2(G155gat), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n860), .B2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n851), .B2(new_n577), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n577), .A2(G162gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n856), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n705), .A2(new_n457), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n452), .B(new_n903), .C1(new_n807), .C2(new_n808), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(new_n506), .ZN(new_n905));
  INV_X1    g704(.A(G169gat), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(new_n268), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n903), .A2(new_n452), .A3(new_n525), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n849), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n667), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n907), .A2(new_n910), .ZN(G1348gat));
  INV_X1    g710(.A(G176gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n904), .A2(new_n912), .A3(new_n768), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n639), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n912), .ZN(G1349gat));
  OAI21_X1  g714(.A(G183gat), .B1(new_n905), .B2(new_n664), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n909), .A2(new_n353), .A3(new_n609), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n506), .A3(new_n577), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n354), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT123), .B(G190gat), .C1(new_n905), .C2(new_n577), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n922), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n849), .A2(new_n354), .A3(new_n576), .A4(new_n908), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT122), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(G1351gat));
  INV_X1    g729(.A(new_n903), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n809), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n853), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n934), .A2(G197gat), .A3(new_n668), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n931), .A2(new_n507), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n889), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n937), .B2(new_n268), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G197gat), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n937), .A2(KEYINPUT125), .A3(new_n268), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  AND2_X1   g740(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n942));
  NOR2_X1   g741(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n934), .A2(G204gat), .A3(new_n665), .ZN(new_n945));
  MUX2_X1   g744(.A(new_n944), .B(new_n942), .S(new_n945), .Z(new_n946));
  OAI21_X1  g745(.A(G204gat), .B1(new_n937), .B2(new_n665), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n889), .A2(new_n609), .A3(new_n936), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n609), .A2(new_n346), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n950), .A2(new_n951), .B1(new_n934), .B2(new_n952), .ZN(G1354gat));
  NAND4_X1  g752(.A1(new_n932), .A2(new_n347), .A3(new_n576), .A4(new_n933), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n889), .A2(new_n955), .A3(new_n936), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n889), .B2(new_n936), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(new_n577), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n958), .B2(new_n347), .ZN(G1355gat));
endmodule


