

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(n754), .ZN(n516) );
  XOR2_X2 U550 ( .A(KEYINPUT17), .B(n517), .Z(n859) );
  XNOR2_X1 U551 ( .A(KEYINPUT32), .B(n763), .ZN(n785) );
  NOR2_X1 U552 ( .A1(n649), .A2(n543), .ZN(n655) );
  NAND2_X1 U553 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U554 ( .A1(n712), .A2(n711), .ZN(n754) );
  INV_X1 U555 ( .A(KEYINPUT98), .ZN(n733) );
  INV_X1 U556 ( .A(KEYINPUT99), .ZN(n737) );
  XNOR2_X1 U557 ( .A(n737), .B(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U558 ( .A(KEYINPUT13), .B(KEYINPUT76), .ZN(n587) );
  XNOR2_X1 U559 ( .A(n588), .B(n587), .ZN(n589) );
  NOR2_X1 U560 ( .A1(n528), .A2(n527), .ZN(G160) );
  AND2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n863) );
  NAND2_X1 U562 ( .A1(G113), .A2(n863), .ZN(n519) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NAND2_X1 U564 ( .A1(G137), .A2(n859), .ZN(n518) );
  NAND2_X1 U565 ( .A1(n519), .A2(n518), .ZN(n528) );
  AND2_X1 U566 ( .A1(G101), .A2(G2104), .ZN(n520) );
  NAND2_X1 U567 ( .A1(n520), .A2(n522), .ZN(n521) );
  XOR2_X1 U568 ( .A(KEYINPUT23), .B(n521), .Z(n524) );
  INV_X1 U569 ( .A(G2105), .ZN(n522) );
  NOR2_X2 U570 ( .A1(G2104), .A2(n522), .ZN(n866) );
  NAND2_X1 U571 ( .A1(n866), .A2(G125), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n526) );
  INV_X1 U573 ( .A(KEYINPUT67), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U575 ( .A(G2427), .B(KEYINPUT104), .ZN(n538) );
  XOR2_X1 U576 ( .A(G2443), .B(G2438), .Z(n530) );
  XNOR2_X1 U577 ( .A(G2430), .B(G2454), .ZN(n529) );
  XNOR2_X1 U578 ( .A(n530), .B(n529), .ZN(n534) );
  XOR2_X1 U579 ( .A(KEYINPUT103), .B(G2435), .Z(n532) );
  XNOR2_X1 U580 ( .A(G1348), .B(G1341), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U582 ( .A(n534), .B(n533), .Z(n536) );
  XNOR2_X1 U583 ( .A(G2451), .B(G2446), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U585 ( .A(n538), .B(n537), .ZN(n539) );
  AND2_X1 U586 ( .A1(n539), .A2(G14), .ZN(G401) );
  INV_X1 U587 ( .A(G651), .ZN(n543) );
  NOR2_X1 U588 ( .A1(G543), .A2(n543), .ZN(n540) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n540), .Z(n656) );
  NAND2_X1 U590 ( .A1(G64), .A2(n656), .ZN(n542) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n649) );
  NOR2_X1 U592 ( .A1(G651), .A2(n649), .ZN(n653) );
  NAND2_X1 U593 ( .A1(G52), .A2(n653), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n549) );
  NAND2_X1 U595 ( .A1(G77), .A2(n655), .ZN(n546) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n544) );
  XNOR2_X1 U597 ( .A(n544), .B(KEYINPUT66), .ZN(n659) );
  NAND2_X1 U598 ( .A1(G90), .A2(n659), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U601 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U603 ( .A1(G111), .A2(n863), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G135), .A2(n859), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n866), .A2(G123), .ZN(n552) );
  XOR2_X1 U607 ( .A(KEYINPUT18), .B(n552), .Z(n553) );
  NOR2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n556) );
  AND2_X1 U609 ( .A1(n522), .A2(G2104), .ZN(n559) );
  NAND2_X1 U610 ( .A1(n559), .A2(G99), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n951) );
  XNOR2_X1 U612 ( .A(G2096), .B(n951), .ZN(n557) );
  OR2_X1 U613 ( .A1(G2100), .A2(n557), .ZN(G156) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  NAND2_X1 U616 ( .A1(G126), .A2(n866), .ZN(n558) );
  XNOR2_X1 U617 ( .A(n558), .B(KEYINPUT86), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G102), .A2(n559), .ZN(n560) );
  XOR2_X1 U619 ( .A(KEYINPUT87), .B(n560), .Z(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n859), .A2(G138), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n863), .A2(G114), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(G164) );
  NAND2_X1 U625 ( .A1(G89), .A2(n659), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U627 ( .A1(G76), .A2(n655), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U629 ( .A(n570), .B(KEYINPUT5), .ZN(n576) );
  XNOR2_X1 U630 ( .A(KEYINPUT6), .B(KEYINPUT79), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G63), .A2(n656), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G51), .A2(n653), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U636 ( .A(KEYINPUT7), .B(n577), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n832) );
  NAND2_X1 U641 ( .A1(n832), .A2(G567), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U643 ( .A1(n656), .A2(G56), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT14), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G43), .A2(n653), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n590) );
  NAND2_X1 U647 ( .A1(n655), .A2(G68), .ZN(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT75), .B(n583), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G81), .A2(n659), .ZN(n584) );
  XOR2_X1 U650 ( .A(n584), .B(KEYINPUT12), .Z(n585) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n588) );
  NOR2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U653 ( .A(KEYINPUT77), .B(n591), .ZN(n988) );
  INV_X1 U654 ( .A(n988), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n592), .A2(G860), .ZN(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G92), .A2(n659), .ZN(n599) );
  NAND2_X1 U659 ( .A1(G66), .A2(n656), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G54), .A2(n653), .ZN(n593) );
  NAND2_X1 U661 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n655), .A2(G79), .ZN(n595) );
  XOR2_X1 U663 ( .A(KEYINPUT78), .B(n595), .Z(n596) );
  NOR2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n600), .Z(n995) );
  INV_X1 U667 ( .A(G868), .ZN(n675) );
  NAND2_X1 U668 ( .A1(n995), .A2(n675), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n656), .A2(G65), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT72), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G53), .A2(n653), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U674 ( .A(KEYINPUT73), .B(n606), .ZN(n611) );
  NAND2_X1 U675 ( .A1(G78), .A2(n655), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G91), .A2(n659), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U678 ( .A(KEYINPUT71), .B(n609), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(G299) );
  NOR2_X1 U680 ( .A1(G286), .A2(n675), .ZN(n613) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U682 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U683 ( .A(G559), .ZN(n616) );
  NOR2_X1 U684 ( .A1(G860), .A2(n616), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n995), .A2(n614), .ZN(n615) );
  XOR2_X1 U686 ( .A(KEYINPUT16), .B(n615), .Z(G148) );
  INV_X1 U687 ( .A(n995), .ZN(n626) );
  NAND2_X1 U688 ( .A1(n616), .A2(n626), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n617), .A2(G868), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n988), .A2(n675), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G67), .A2(n656), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G55), .A2(n653), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U695 ( .A1(G80), .A2(n655), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G93), .A2(n659), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n674) );
  NAND2_X1 U699 ( .A1(G559), .A2(n626), .ZN(n627) );
  XOR2_X1 U700 ( .A(n988), .B(n627), .Z(n672) );
  XOR2_X1 U701 ( .A(n672), .B(KEYINPUT80), .Z(n628) );
  NOR2_X1 U702 ( .A1(G860), .A2(n628), .ZN(n629) );
  XOR2_X1 U703 ( .A(n674), .B(n629), .Z(G145) );
  NAND2_X1 U704 ( .A1(G72), .A2(n655), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G85), .A2(n659), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n637) );
  NAND2_X1 U707 ( .A1(n653), .A2(G47), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT68), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G60), .A2(n656), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT69), .B(n635), .Z(n636) );
  NOR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U713 ( .A(KEYINPUT70), .B(n638), .Z(G290) );
  NAND2_X1 U714 ( .A1(G61), .A2(n656), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G48), .A2(n653), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n655), .A2(G73), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G86), .A2(n659), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G49), .A2(n653), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U725 ( .A1(n656), .A2(n648), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G87), .A2(n649), .ZN(n650) );
  XOR2_X1 U727 ( .A(KEYINPUT81), .B(n650), .Z(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G50), .A2(n653), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(KEYINPUT82), .ZN(n664) );
  NAND2_X1 U731 ( .A1(G75), .A2(n655), .ZN(n658) );
  NAND2_X1 U732 ( .A1(G62), .A2(n656), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U734 ( .A1(G88), .A2(n659), .ZN(n660) );
  XNOR2_X1 U735 ( .A(KEYINPUT83), .B(n660), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT84), .B(n665), .ZN(G303) );
  XOR2_X1 U739 ( .A(n674), .B(G305), .Z(n668) );
  XNOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n666), .B(G288), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U743 ( .A(G290), .B(n669), .ZN(n671) );
  XNOR2_X1 U744 ( .A(G299), .B(G303), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(n882) );
  XNOR2_X1 U746 ( .A(n672), .B(n882), .ZN(n673) );
  NAND2_X1 U747 ( .A1(n673), .A2(G868), .ZN(n677) );
  NAND2_X1 U748 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U749 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U754 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U756 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U759 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U760 ( .A1(G96), .A2(n684), .ZN(n836) );
  NAND2_X1 U761 ( .A1(n836), .A2(G2106), .ZN(n688) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U763 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U764 ( .A1(G108), .A2(n686), .ZN(n837) );
  NAND2_X1 U765 ( .A1(n837), .A2(G567), .ZN(n687) );
  NAND2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n886) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U768 ( .A1(n886), .A2(n689), .ZN(n835) );
  NAND2_X1 U769 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G107), .A2(n863), .ZN(n691) );
  NAND2_X1 U771 ( .A1(G119), .A2(n866), .ZN(n690) );
  NAND2_X1 U772 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U773 ( .A(KEYINPUT91), .B(n692), .ZN(n697) );
  NAND2_X1 U774 ( .A1(G95), .A2(n559), .ZN(n694) );
  NAND2_X1 U775 ( .A1(G131), .A2(n859), .ZN(n693) );
  NAND2_X1 U776 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U777 ( .A(KEYINPUT92), .B(n695), .Z(n696) );
  NAND2_X1 U778 ( .A1(n697), .A2(n696), .ZN(n873) );
  NAND2_X1 U779 ( .A1(G1991), .A2(n873), .ZN(n698) );
  XNOR2_X1 U780 ( .A(KEYINPUT93), .B(n698), .ZN(n708) );
  NAND2_X1 U781 ( .A1(G117), .A2(n863), .ZN(n700) );
  NAND2_X1 U782 ( .A1(G141), .A2(n859), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U784 ( .A1(n559), .A2(G105), .ZN(n701) );
  XOR2_X1 U785 ( .A(KEYINPUT38), .B(n701), .Z(n702) );
  NOR2_X1 U786 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U787 ( .A1(n866), .A2(G129), .ZN(n704) );
  NAND2_X1 U788 ( .A1(n705), .A2(n704), .ZN(n874) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n874), .ZN(n706) );
  XOR2_X1 U790 ( .A(KEYINPUT94), .B(n706), .Z(n707) );
  NOR2_X1 U791 ( .A1(n708), .A2(n707), .ZN(n943) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NAND2_X1 U793 ( .A1(G160), .A2(G40), .ZN(n709) );
  NOR2_X1 U794 ( .A1(n711), .A2(n709), .ZN(n823) );
  INV_X1 U795 ( .A(n823), .ZN(n710) );
  NOR2_X1 U796 ( .A1(n943), .A2(n710), .ZN(n818) );
  AND2_X1 U797 ( .A1(G160), .A2(G40), .ZN(n712) );
  NAND2_X1 U798 ( .A1(n516), .A2(G2072), .ZN(n713) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(n713), .Z(n715) );
  NAND2_X1 U800 ( .A1(G1956), .A2(n754), .ZN(n714) );
  NAND2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n728) );
  NAND2_X1 U802 ( .A1(G299), .A2(n728), .ZN(n716) );
  XOR2_X1 U803 ( .A(KEYINPUT28), .B(n716), .Z(n736) );
  NAND2_X1 U804 ( .A1(n516), .A2(G1996), .ZN(n718) );
  XOR2_X1 U805 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n717) );
  XNOR2_X1 U806 ( .A(n718), .B(n717), .ZN(n720) );
  NAND2_X1 U807 ( .A1(n754), .A2(G1341), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U809 ( .A(KEYINPUT97), .B(n721), .Z(n722) );
  NOR2_X1 U810 ( .A1(n988), .A2(n722), .ZN(n726) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n754), .ZN(n724) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n516), .ZN(n723) );
  NAND2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U814 ( .A1(n995), .A2(n727), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n732) );
  NOR2_X1 U816 ( .A1(n995), .A2(n727), .ZN(n730) );
  NOR2_X1 U817 ( .A1(n728), .A2(G299), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U819 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n739) );
  XNOR2_X1 U821 ( .A(n739), .B(n738), .ZN(n745) );
  NOR2_X1 U822 ( .A1(n516), .A2(G1961), .ZN(n740) );
  XNOR2_X1 U823 ( .A(n740), .B(KEYINPUT95), .ZN(n743) );
  XNOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .ZN(n741) );
  XNOR2_X1 U825 ( .A(n741), .B(KEYINPUT96), .ZN(n915) );
  NAND2_X1 U826 ( .A1(n915), .A2(n516), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n743), .A2(n742), .ZN(n749) );
  NAND2_X1 U828 ( .A1(G171), .A2(n749), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n765) );
  NAND2_X1 U830 ( .A1(G8), .A2(n754), .ZN(n793) );
  NOR2_X1 U831 ( .A1(G1966), .A2(n793), .ZN(n767) );
  NOR2_X1 U832 ( .A1(G2084), .A2(n754), .ZN(n766) );
  NOR2_X1 U833 ( .A1(n767), .A2(n766), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U835 ( .A(KEYINPUT30), .B(n747), .ZN(n748) );
  NOR2_X1 U836 ( .A1(G168), .A2(n748), .ZN(n751) );
  NOR2_X1 U837 ( .A1(G171), .A2(n749), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U839 ( .A(KEYINPUT31), .B(n752), .Z(n764) );
  NAND2_X1 U840 ( .A1(n765), .A2(n764), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n753), .A2(G286), .ZN(n762) );
  INV_X1 U842 ( .A(G8), .ZN(n760) );
  NOR2_X1 U843 ( .A1(G2090), .A2(n754), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(KEYINPUT100), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n793), .A2(G1971), .ZN(n756) );
  NOR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n758), .A2(G303), .ZN(n759) );
  OR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U850 ( .A1(n765), .A2(n764), .ZN(n770) );
  AND2_X1 U851 ( .A1(G8), .A2(n766), .ZN(n768) );
  OR2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U853 ( .A1(n770), .A2(n769), .ZN(n786) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n998) );
  INV_X1 U855 ( .A(n793), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n998), .A2(n771), .ZN(n775) );
  INV_X1 U857 ( .A(n775), .ZN(n772) );
  AND2_X1 U858 ( .A1(n786), .A2(n772), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n785), .A2(n773), .ZN(n777) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n780) );
  NOR2_X1 U861 ( .A1(G303), .A2(G1971), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n780), .A2(n774), .ZN(n1004) );
  OR2_X1 U863 ( .A1(n775), .A2(n1004), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n778), .B(KEYINPUT64), .ZN(n779) );
  NOR2_X1 U866 ( .A1(KEYINPUT33), .A2(n779), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n780), .A2(KEYINPUT33), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n781), .A2(n793), .ZN(n782) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U870 ( .A(G1981), .B(G305), .Z(n989) );
  AND2_X1 U871 ( .A1(n784), .A2(n989), .ZN(n797) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G8), .A2(n787), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U876 ( .A1(n790), .A2(n793), .ZN(n795) );
  NOR2_X1 U877 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XOR2_X1 U878 ( .A(n791), .B(KEYINPUT24), .Z(n792) );
  OR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U882 ( .A1(n818), .A2(n798), .ZN(n813) );
  XNOR2_X1 U883 ( .A(KEYINPUT88), .B(G290), .ZN(n799) );
  XNOR2_X1 U884 ( .A(n799), .B(G1986), .ZN(n1010) );
  NAND2_X1 U885 ( .A1(n1010), .A2(n823), .ZN(n811) );
  NAND2_X1 U886 ( .A1(G116), .A2(n863), .ZN(n801) );
  NAND2_X1 U887 ( .A1(G128), .A2(n866), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n802), .Z(n809) );
  NAND2_X1 U890 ( .A1(G140), .A2(n859), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n559), .A2(G104), .ZN(n803) );
  XOR2_X1 U892 ( .A(KEYINPUT89), .B(n803), .Z(n804) );
  NAND2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(KEYINPUT34), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(KEYINPUT90), .ZN(n808) );
  NOR2_X1 U896 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U897 ( .A(KEYINPUT36), .B(n810), .Z(n877) );
  XOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .Z(n822) );
  AND2_X1 U899 ( .A1(n877), .A2(n822), .ZN(n940) );
  NAND2_X1 U900 ( .A1(n940), .A2(n823), .ZN(n814) );
  AND2_X1 U901 ( .A1(n811), .A2(n814), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n829) );
  INV_X1 U903 ( .A(n814), .ZN(n827) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n874), .ZN(n947) );
  NOR2_X1 U905 ( .A1(G290), .A2(G1986), .ZN(n815) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n873), .ZN(n953) );
  NOR2_X1 U907 ( .A1(n815), .A2(n953), .ZN(n816) );
  XOR2_X1 U908 ( .A(KEYINPUT101), .B(n816), .Z(n817) );
  NOR2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U910 ( .A1(n947), .A2(n819), .ZN(n820) );
  XNOR2_X1 U911 ( .A(KEYINPUT39), .B(n820), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n821), .A2(n823), .ZN(n825) );
  NOR2_X1 U913 ( .A1(n877), .A2(n822), .ZN(n941) );
  NAND2_X1 U914 ( .A1(n941), .A2(n823), .ZN(n824) );
  AND2_X1 U915 ( .A1(n825), .A2(n824), .ZN(n826) );
  OR2_X1 U916 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n829), .A2(n828), .ZN(n831) );
  XNOR2_X1 U918 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n830) );
  XNOR2_X1 U919 ( .A(n831), .B(n830), .ZN(G329) );
  INV_X1 U920 ( .A(G303), .ZN(G166) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U923 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U925 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  NAND2_X1 U932 ( .A1(G124), .A2(n866), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT105), .B(n838), .Z(n839) );
  XNOR2_X1 U934 ( .A(n839), .B(KEYINPUT44), .ZN(n841) );
  NAND2_X1 U935 ( .A1(G112), .A2(n863), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U937 ( .A1(G100), .A2(n559), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G136), .A2(n859), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G162) );
  XOR2_X1 U941 ( .A(G160), .B(G162), .Z(n846) );
  XNOR2_X1 U942 ( .A(n951), .B(n846), .ZN(n850) );
  XOR2_X1 U943 ( .A(KEYINPUT48), .B(KEYINPUT107), .Z(n848) );
  XNOR2_X1 U944 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(n850), .B(n849), .Z(n872) );
  NAND2_X1 U947 ( .A1(G103), .A2(n559), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G139), .A2(n859), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U950 ( .A1(G115), .A2(n863), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G127), .A2(n866), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(KEYINPUT47), .B(n855), .Z(n856) );
  NOR2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U955 ( .A(KEYINPUT109), .B(n858), .Z(n935) );
  NAND2_X1 U956 ( .A1(G106), .A2(n559), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G142), .A2(n859), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n862), .B(KEYINPUT45), .ZN(n865) );
  NAND2_X1 U960 ( .A1(G118), .A2(n863), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U962 ( .A1(n866), .A2(G130), .ZN(n867) );
  XOR2_X1 U963 ( .A(KEYINPUT106), .B(n867), .Z(n868) );
  NOR2_X1 U964 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U965 ( .A(n935), .B(n870), .ZN(n871) );
  XNOR2_X1 U966 ( .A(n872), .B(n871), .ZN(n879) );
  XNOR2_X1 U967 ( .A(G164), .B(n873), .ZN(n875) );
  XNOR2_X1 U968 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U969 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U970 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U971 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U972 ( .A(G286), .B(n995), .ZN(n881) );
  XNOR2_X1 U973 ( .A(n881), .B(G301), .ZN(n884) );
  XNOR2_X1 U974 ( .A(n988), .B(n882), .ZN(n883) );
  XNOR2_X1 U975 ( .A(n884), .B(n883), .ZN(n885) );
  NOR2_X1 U976 ( .A1(G37), .A2(n885), .ZN(G397) );
  INV_X1 U977 ( .A(n886), .ZN(G319) );
  XOR2_X1 U978 ( .A(G2100), .B(G2096), .Z(n888) );
  XNOR2_X1 U979 ( .A(KEYINPUT42), .B(G2678), .ZN(n887) );
  XNOR2_X1 U980 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U981 ( .A(KEYINPUT43), .B(G2090), .Z(n890) );
  XNOR2_X1 U982 ( .A(G2067), .B(G2072), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U984 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U985 ( .A(G2078), .B(G2084), .ZN(n893) );
  XNOR2_X1 U986 ( .A(n894), .B(n893), .ZN(G227) );
  XOR2_X1 U987 ( .A(G1986), .B(G1976), .Z(n896) );
  XNOR2_X1 U988 ( .A(G1956), .B(G1971), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U990 ( .A(n897), .B(G2474), .Z(n899) );
  XNOR2_X1 U991 ( .A(G1966), .B(G1981), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U993 ( .A(KEYINPUT41), .B(G1991), .Z(n901) );
  XNOR2_X1 U994 ( .A(G1996), .B(G1961), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(G229) );
  NOR2_X1 U997 ( .A1(G395), .A2(G397), .ZN(n904) );
  XOR2_X1 U998 ( .A(KEYINPUT111), .B(n904), .Z(n910) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n905) );
  XOR2_X1 U1000 ( .A(KEYINPUT49), .B(n905), .Z(n906) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n906), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(KEYINPUT110), .B(n908), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1007 ( .A(KEYINPUT55), .B(KEYINPUT114), .Z(n959) );
  XNOR2_X1 U1008 ( .A(KEYINPUT115), .B(G2090), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(G35), .ZN(n928) );
  XOR2_X1 U1010 ( .A(G1991), .B(KEYINPUT116), .Z(n912) );
  XNOR2_X1 U1011 ( .A(G25), .B(n912), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n913), .A2(G28), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n914), .B(KEYINPUT117), .ZN(n924) );
  XNOR2_X1 U1014 ( .A(n915), .B(G27), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(G2072), .B(G33), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G32), .B(G1996), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT118), .B(G2067), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(G26), .B(n920), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n925) );
  XNOR2_X1 U1024 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(G34), .B(G2084), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT54), .B(n929), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n959), .B(n932), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(G29), .A2(n933), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT120), .B(n934), .Z(n963) );
  XNOR2_X1 U1032 ( .A(G2072), .B(n935), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(G164), .B(G2078), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n936), .B(KEYINPUT112), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(n939), .B(KEYINPUT50), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n956) );
  XOR2_X1 U1040 ( .A(G160), .B(G2084), .Z(n950) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT51), .B(n948), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n954) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n957), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n958), .B(KEYINPUT113), .ZN(n960) );
  NAND2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1051 ( .A1(n961), .A2(G29), .ZN(n962) );
  NAND2_X1 U1052 ( .A1(n963), .A2(n962), .ZN(n1018) );
  XOR2_X1 U1053 ( .A(G1348), .B(KEYINPUT59), .Z(n964) );
  XNOR2_X1 U1054 ( .A(G4), .B(n964), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G20), .B(G1956), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n970) );
  XNOR2_X1 U1057 ( .A(G1341), .B(G19), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G1981), .B(G6), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n971), .B(KEYINPUT60), .ZN(n985) );
  XOR2_X1 U1062 ( .A(G1986), .B(G24), .Z(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(n972), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(G1976), .B(G23), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT124), .B(n975), .Z(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(KEYINPUT126), .B(n978), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n979), .B(KEYINPUT58), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G5), .B(G1961), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1076 ( .A(KEYINPUT61), .B(n986), .Z(n987) );
  NOR2_X1 U1077 ( .A1(G16), .A2(n987), .ZN(n1015) );
  XOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .Z(n1012) );
  XNOR2_X1 U1079 ( .A(n988), .B(G1341), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n991), .B(KEYINPUT121), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT57), .B(n992), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n1008) );
  NAND2_X1 U1085 ( .A1(G303), .A2(G1971), .ZN(n997) );
  XOR2_X1 U1086 ( .A(G1348), .B(n995), .Z(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G171), .B(G1961), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G299), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(KEYINPUT122), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(KEYINPUT123), .B(n1013), .Z(n1014) );
  NOR2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(n1016), .B(KEYINPUT127), .ZN(n1017) );
  NOR2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(G11), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

