//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n455), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n463), .B2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n467), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(new_n471), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n484), .A3(new_n471), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(new_n471), .B2(G112), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n487), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT71), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n471), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n500), .B1(new_n482), .B2(G126), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n501), .B2(new_n471), .ZN(new_n502));
  OAI21_X1  g077(.A(G138), .B1(KEYINPUT72), .B2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n482), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(G102), .A2(G2104), .ZN(new_n507));
  AOI21_X1  g082(.A(G2105), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n502), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(G651), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n513), .A2(KEYINPUT74), .A3(KEYINPUT6), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(new_n511), .B2(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(G543), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  OAI21_X1  g099(.A(G543), .B1(new_n524), .B2(KEYINPUT75), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(new_n515), .A3(new_n519), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G62), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n522), .B1(new_n523), .B2(new_n531), .C1(new_n536), .C2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND3_X1  g114(.A1(new_n515), .A2(G89), .A3(new_n519), .ZN(new_n540));
  INV_X1    g115(.A(G63), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n513), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(new_n530), .B1(new_n521), .B2(G51), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G168));
  INV_X1    g123(.A(new_n531), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(G90), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n529), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(G171));
  NAND2_X1  g133(.A1(new_n549), .A2(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n521), .A2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n529), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n529), .B(KEYINPUT79), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G91), .B2(new_n549), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n520), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n557), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT80), .A4(new_n556), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G301));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n547), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n543), .A2(KEYINPUT81), .A3(new_n546), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G286));
  OAI21_X1  g165(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n530), .A2(new_n515), .A3(G87), .A4(new_n519), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n515), .A2(G49), .A3(G543), .A4(new_n519), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  NAND3_X1  g169(.A1(new_n515), .A2(G48), .A3(new_n519), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G651), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n527), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n515), .A2(G86), .A3(new_n519), .ZN(new_n598));
  NAND2_X1  g173(.A1(G61), .A2(G651), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n529), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n549), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n521), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n529), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n603), .A2(new_n604), .A3(new_n608), .ZN(G290));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  NOR3_X1   g186(.A1(new_n531), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n610), .B1(new_n531), .B2(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n521), .A2(G54), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n574), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G651), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n615), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G301), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G284));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(new_n622), .ZN(G321));
  MUX2_X1   g201(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g202(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g203(.A(new_n621), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g210(.A(new_n486), .ZN(new_n636));
  INV_X1    g211(.A(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(KEYINPUT85), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n486), .A2(new_n639), .A3(G123), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n638), .A2(new_n640), .B1(G135), .B2(new_n489), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n642));
  OR2_X1    g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n641), .B2(new_n644), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n473), .A2(new_n482), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT13), .Z(new_n652));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n653), .A2(G2100), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(G2100), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n648), .B(new_n656), .C1(new_n654), .C2(new_n652), .ZN(G156));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT87), .B(G2438), .Z(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT15), .B(G2435), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT14), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(G14), .ZN(G401));
  XOR2_X1   g246(.A(G2067), .B(G2678), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(KEYINPUT17), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(new_n675), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n676), .B(KEYINPUT88), .Z(new_n683));
  OAI211_X1 g258(.A(new_n678), .B(new_n682), .C1(new_n680), .C2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(new_n688), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n688), .A3(new_n691), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G19), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n566), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G1341), .ZN(new_n710));
  AND2_X1   g285(.A1(KEYINPUT91), .A2(G29), .ZN(new_n711));
  NOR2_X1   g286(.A1(KEYINPUT91), .A2(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT29), .Z(new_n717));
  INV_X1    g292(.A(G2090), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n714), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT100), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2078), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT98), .B(G34), .Z(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT24), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT24), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n725), .A2(new_n714), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n479), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G2084), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G28), .ZN(new_n732));
  AOI21_X1  g307(.A(G29), .B1(new_n732), .B2(KEYINPUT30), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(KEYINPUT30), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n730), .B2(new_n729), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT31), .B(G11), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n739));
  INV_X1    g314(.A(G26), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n713), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n714), .A2(KEYINPUT28), .A3(G26), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n486), .A2(G128), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n489), .A2(G140), .ZN(new_n744));
  OR2_X1    g319(.A1(G104), .A2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n741), .B(new_n742), .C1(new_n748), .C2(new_n728), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n728), .A2(G33), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT25), .Z(new_n753));
  AOI22_X1  g328(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  INV_X1    g329(.A(G139), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n753), .B1(new_n471), .B2(new_n754), .C1(new_n488), .C2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(new_n728), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n750), .B1(G2072), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n647), .A2(new_n713), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n737), .A2(new_n738), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n486), .A2(G129), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n489), .A2(G141), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n473), .A2(G105), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n764), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G29), .B2(G32), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT27), .B(G1996), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT99), .ZN(new_n774));
  NAND2_X1  g349(.A1(G171), .A2(G16), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G5), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n772), .A2(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G21), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G168), .B2(G16), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n772), .A2(new_n774), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n780), .A2(G1966), .B1(new_n709), .B2(G1341), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n776), .A2(new_n777), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n763), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n707), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n629), .B2(new_n707), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1348), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n707), .A2(G20), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT101), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT23), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n760), .A2(KEYINPUT97), .A3(G2072), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT97), .B1(new_n760), .B2(G2072), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n790), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n717), .A2(new_n718), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n719), .A2(new_n787), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n802));
  INV_X1    g377(.A(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G16), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G303), .B2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n804), .B1(new_n806), .B2(new_n802), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G1971), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n707), .A2(G6), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n601), .B2(new_n707), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT32), .B(G1981), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n807), .A2(G1971), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT93), .B1(G16), .B2(G23), .ZN(new_n814));
  OR3_X1    g389(.A1(KEYINPUT93), .A2(G16), .A3(G23), .ZN(new_n815));
  NAND2_X1  g390(.A1(G288), .A2(KEYINPUT94), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n817), .A4(new_n593), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n814), .B(new_n815), .C1(new_n820), .C2(new_n707), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT33), .B(G1976), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n808), .A2(new_n812), .A3(new_n813), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  AOI22_X1  g400(.A1(G119), .A2(new_n486), .B1(new_n489), .B2(G131), .ZN(new_n826));
  OR2_X1    g401(.A1(G95), .A2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT92), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G25), .B(new_n830), .S(new_n713), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT35), .B(G1991), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n707), .A2(G24), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n707), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(G1986), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G1986), .B2(new_n836), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n824), .B2(KEYINPUT34), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n831), .A2(new_n832), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n825), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n843));
  AOI211_X1 g418(.A(new_n710), .B(new_n801), .C1(new_n842), .C2(new_n843), .ZN(G311));
  AOI21_X1  g419(.A(new_n801), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G1341), .B2(new_n709), .ZN(G150));
  XNOR2_X1  g421(.A(KEYINPUT102), .B(G93), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n549), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n521), .A2(G55), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n848), .B(new_n849), .C1(new_n513), .C2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT103), .B(G860), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n565), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n621), .A2(new_n630), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n854), .B1(new_n859), .B2(new_n852), .ZN(G145));
  NAND2_X1  g435(.A1(new_n486), .A2(G130), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n489), .A2(G142), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n471), .A2(G118), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n463), .B1(new_n863), .B2(KEYINPUT105), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n864), .B1(KEYINPUT105), .B2(new_n863), .C1(G106), .C2(G2105), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n651), .ZN(new_n867));
  OAI21_X1  g442(.A(G160), .B1(new_n645), .B2(new_n646), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT86), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n479), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n769), .B(new_n747), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT104), .B1(new_n502), .B2(new_n508), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n499), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n876), .A2(G2105), .B1(new_n497), .B2(new_n496), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n464), .A2(new_n466), .A3(new_n505), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n507), .B1(new_n878), .B2(new_n503), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n471), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n873), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n874), .A2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n770), .A2(new_n747), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n748), .A2(new_n769), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n883), .A2(new_n756), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n758), .B1(new_n883), .B2(new_n887), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n868), .B(new_n872), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n883), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n759), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n868), .A2(new_n872), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n883), .A2(new_n887), .A3(new_n756), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n494), .B(new_n830), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n890), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n890), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n867), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n896), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n867), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n890), .A2(new_n895), .A3(new_n896), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n899), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n621), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n613), .A2(new_n614), .B1(new_n619), .B2(G651), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(new_n581), .A3(new_n577), .A4(new_n616), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n911), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n911), .A2(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT106), .B1(new_n918), .B2(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n632), .B(new_n855), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n918), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OR3_X1    g499(.A1(new_n922), .A2(KEYINPUT42), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n835), .A2(G305), .ZN(new_n926));
  NAND2_X1  g501(.A1(G290), .A2(new_n601), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n819), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n819), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(G303), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(G166), .A3(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n922), .B2(new_n924), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n925), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n925), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n851), .A2(new_n622), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  INV_X1    g517(.A(new_n589), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT81), .B1(new_n543), .B2(new_n546), .ZN(new_n944));
  OAI21_X1  g519(.A(G171), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n547), .B1(new_n584), .B2(new_n585), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n947), .A3(new_n855), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n566), .B(new_n851), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n557), .B1(new_n588), .B2(new_n589), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(new_n946), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n917), .A2(new_n919), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n918), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n948), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n934), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n948), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT106), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n919), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n934), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n963), .A3(new_n954), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n956), .A2(new_n907), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n958), .A2(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n957), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(KEYINPUT107), .A3(new_n954), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n951), .A2(new_n948), .A3(new_n953), .A4(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n934), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(new_n964), .A3(new_n907), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n942), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n942), .B1(new_n975), .B2(KEYINPUT43), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n956), .A2(new_n964), .A3(new_n966), .A4(new_n907), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n978), .A2(KEYINPUT108), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT108), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(G397));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n884), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT109), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n474), .A2(G40), .A3(new_n478), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n884), .A2(new_n989), .A3(new_n983), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n985), .A2(new_n986), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G2067), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n747), .B(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT110), .ZN(new_n995));
  INV_X1    g570(.A(new_n991), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n830), .A2(new_n832), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n830), .A2(new_n832), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n769), .B(G1996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(G290), .B(G1986), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n996), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n577), .A2(new_n1005), .A3(new_n581), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n577), .B2(new_n581), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n877), .B2(new_n880), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n983), .B1(new_n502), .B2(new_n508), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1013), .A3(new_n988), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n795), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n502), .A2(new_n508), .A3(KEYINPUT104), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n881), .B1(new_n877), .B2(new_n880), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT45), .B(new_n983), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n884), .A2(new_n1020), .A3(KEYINPUT45), .A4(new_n983), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1012), .A2(KEYINPUT111), .A3(new_n986), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1019), .A2(new_n988), .A3(new_n1021), .A4(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1008), .B(new_n1015), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1015), .ZN(new_n1030));
  AND4_X1   g605(.A1(new_n988), .A2(new_n1019), .A3(new_n1021), .A4(new_n1025), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n1027), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(new_n1008), .ZN(new_n1033));
  INV_X1    g608(.A(G1348), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1012), .A2(new_n987), .A3(G2067), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1014), .A2(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1036), .A2(new_n1035), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n621), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1029), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(KEYINPUT60), .A3(new_n1038), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT60), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n621), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(KEYINPUT60), .A3(new_n629), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT119), .B(G1996), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1012), .A2(new_n987), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT58), .B(G1341), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1026), .A2(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n566), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1050), .B2(new_n566), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1046), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT61), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1032), .A2(KEYINPUT120), .A3(new_n1055), .A4(new_n1008), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT61), .B1(new_n1029), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1041), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT113), .B(G1971), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1026), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1014), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n718), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G303), .A2(G8), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1066), .B(KEYINPUT55), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1026), .A2(new_n1061), .B1(new_n718), .B2(new_n1063), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT114), .B(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n819), .A2(G1976), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1048), .A2(new_n1073), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT115), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  NAND3_X1  g657(.A1(G288), .A2(new_n1077), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT49), .ZN(new_n1084));
  OAI21_X1  g659(.A(G1981), .B1(new_n597), .B2(new_n600), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n597), .A2(new_n600), .A3(G1981), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1981), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n601), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(KEYINPUT49), .A3(new_n1085), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1091), .A3(new_n1076), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1091), .A3(KEYINPUT116), .A4(new_n1076), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1081), .A2(new_n1083), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1069), .A2(new_n1074), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1012), .A2(new_n986), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT45), .B(new_n983), .C1(new_n502), .C2(new_n508), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n988), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1966), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1011), .A2(new_n1013), .A3(new_n730), .A4(new_n988), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1073), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n547), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1104), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G168), .A2(new_n1073), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1113), .B2(new_n1109), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1104), .A2(KEYINPUT51), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1109), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1097), .B1(new_n1105), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1026), .B2(G2078), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(G2078), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1098), .A2(new_n988), .A3(new_n1099), .A4(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT122), .B(G1961), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1014), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n624), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n985), .A2(new_n986), .A3(new_n990), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n988), .A3(new_n1131), .A4(new_n1124), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1132), .A2(new_n1123), .A3(G301), .A4(new_n1127), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1121), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g711(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1060), .B(new_n1120), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .A3(G301), .A4(new_n1125), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1132), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1135), .B1(new_n1141), .B2(G171), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1128), .B2(new_n624), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT125), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1138), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1117), .B1(new_n1116), .B2(new_n1109), .ZN(new_n1151));
  NOR4_X1   g726(.A1(new_n1104), .A2(KEYINPUT121), .A3(new_n1108), .A4(KEYINPUT51), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1151), .A2(new_n1114), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1105), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT62), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1097), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1129), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1119), .A2(new_n1158), .A3(new_n1105), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1161), .A2(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(KEYINPUT117), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1104), .A2(new_n588), .A3(new_n589), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1162), .B(new_n1163), .C1(new_n1097), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1065), .A2(G8), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1161), .B1(new_n1166), .B2(new_n1070), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1164), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n1069), .A3(new_n1096), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1096), .A2(G8), .A3(new_n1068), .A4(new_n1065), .ZN(new_n1171));
  AOI211_X1 g746(.A(G1976), .B(G288), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1076), .B1(new_n1172), .B2(new_n1087), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1160), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1004), .B1(new_n1150), .B2(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n996), .A2(KEYINPUT48), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT48), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1177), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n991), .B2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n995), .A2(new_n997), .A3(new_n1001), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n747), .A2(G2067), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n996), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT46), .ZN(new_n1187));
  OR3_X1    g762(.A1(new_n991), .A2(new_n1187), .A3(G1996), .ZN(new_n1188));
  INV_X1    g763(.A(new_n993), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n996), .B1(new_n769), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1187), .B1(new_n991), .B2(G1996), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1193));
  XNOR2_X1  g768(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1183), .A2(new_n1186), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1175), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g771(.A1(new_n967), .A2(new_n976), .ZN(new_n1198));
  NOR2_X1   g772(.A1(G401), .A2(G227), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n908), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g774(.A1(G229), .A2(new_n461), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  NOR3_X1   g776(.A1(new_n1198), .A2(new_n1200), .A3(new_n1202), .ZN(G308));
  INV_X1    g777(.A(new_n976), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1204), .B1(new_n966), .B2(new_n965), .ZN(new_n1205));
  NAND4_X1  g779(.A1(new_n1205), .A2(new_n908), .A3(new_n1201), .A4(new_n1199), .ZN(G225));
endmodule


