

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  NOR2_X1 U324 ( .A1(n562), .A2(n590), .ZN(n452) );
  NOR2_X1 U325 ( .A1(n475), .A2(n533), .ZN(n384) );
  XOR2_X1 U326 ( .A(n559), .B(KEYINPUT36), .Z(n590) );
  INV_X1 U327 ( .A(n579), .ZN(n480) );
  INV_X1 U328 ( .A(n591), .ZN(n587) );
  NOR2_X1 U329 ( .A1(n567), .A2(n480), .ZN(n481) );
  XNOR2_X1 U330 ( .A(n395), .B(n394), .ZN(n486) );
  XOR2_X2 U331 ( .A(n472), .B(KEYINPUT28), .Z(n530) );
  XOR2_X1 U332 ( .A(G106GAT), .B(G78GAT), .Z(n437) );
  XNOR2_X1 U333 ( .A(n295), .B(n294), .ZN(n360) );
  INV_X1 U334 ( .A(G197GAT), .ZN(n292) );
  INV_X1 U335 ( .A(KEYINPUT110), .ZN(n465) );
  XNOR2_X1 U336 ( .A(n298), .B(G22GAT), .ZN(n299) );
  XNOR2_X1 U337 ( .A(n465), .B(KEYINPUT48), .ZN(n466) );
  INV_X1 U338 ( .A(KEYINPUT92), .ZN(n394) );
  XNOR2_X1 U339 ( .A(n360), .B(n299), .ZN(n304) );
  XNOR2_X1 U340 ( .A(n467), .B(n466), .ZN(n548) );
  XNOR2_X1 U341 ( .A(n520), .B(KEYINPUT102), .ZN(n529) );
  NOR2_X1 U342 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U343 ( .A(KEYINPUT38), .B(n448), .ZN(n504) );
  XNOR2_X1 U344 ( .A(n477), .B(G176GAT), .ZN(n478) );
  XNOR2_X1 U345 ( .A(n449), .B(KEYINPUT100), .ZN(n450) );
  XNOR2_X1 U346 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  XNOR2_X1 U347 ( .A(n451), .B(n450), .ZN(G1331GAT) );
  XNOR2_X1 U348 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n293), .B(n292), .ZN(n295) );
  XOR2_X1 U350 ( .A(G211GAT), .B(G218GAT), .Z(n294) );
  XOR2_X1 U351 ( .A(KEYINPUT81), .B(KEYINPUT23), .Z(n297) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n301) );
  XOR2_X1 U355 ( .A(G50GAT), .B(G162GAT), .Z(n315) );
  XNOR2_X1 U356 ( .A(n315), .B(n437), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(n302), .B(G148GAT), .Z(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U360 ( .A(KEYINPUT3), .B(KEYINPUT82), .Z(n306) );
  XNOR2_X1 U361 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(n307), .ZN(n379) );
  XNOR2_X1 U364 ( .A(n379), .B(KEYINPUT24), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n472) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .Z(n358) );
  INV_X1 U367 ( .A(G85GAT), .ZN(n310) );
  NAND2_X1 U368 ( .A1(G99GAT), .A2(n310), .ZN(n313) );
  INV_X1 U369 ( .A(G99GAT), .ZN(n311) );
  NAND2_X1 U370 ( .A1(n311), .A2(G85GAT), .ZN(n312) );
  NAND2_X1 U371 ( .A1(n313), .A2(n312), .ZN(n443) );
  XNOR2_X1 U372 ( .A(n358), .B(n443), .ZN(n317) );
  AND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n325) );
  XOR2_X1 U376 ( .A(KEYINPUT10), .B(G92GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(G106GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U379 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n321) );
  XNOR2_X1 U380 ( .A(KEYINPUT65), .B(KEYINPUT67), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U382 ( .A(n323), .B(n322), .Z(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U384 ( .A(KEYINPUT75), .B(KEYINPUT73), .Z(n327) );
  XNOR2_X1 U385 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n326) );
  XOR2_X1 U386 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n333) );
  XNOR2_X1 U388 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n330), .B(KEYINPUT7), .ZN(n423) );
  XNOR2_X1 U390 ( .A(G29GAT), .B(G134GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n331), .B(KEYINPUT74), .ZN(n364) );
  XOR2_X1 U392 ( .A(n423), .B(n364), .Z(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n559) );
  XOR2_X1 U394 ( .A(G15GAT), .B(G71GAT), .Z(n335) );
  NAND2_X1 U395 ( .A1(G227GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U397 ( .A(G176GAT), .B(KEYINPUT64), .Z(n337) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(KEYINPUT20), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U400 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U401 ( .A(G134GAT), .B(G190GAT), .Z(n341) );
  XNOR2_X1 U402 ( .A(G43GAT), .B(G99GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(n342), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n350) );
  XOR2_X1 U406 ( .A(G183GAT), .B(KEYINPUT17), .Z(n346) );
  XNOR2_X1 U407 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n355) );
  XOR2_X1 U409 ( .A(G127GAT), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X1 U410 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n374) );
  XOR2_X1 U412 ( .A(n355), .B(n374), .Z(n349) );
  XOR2_X1 U413 ( .A(n350), .B(n349), .Z(n534) );
  INV_X1 U414 ( .A(n534), .ZN(n475) );
  XOR2_X1 U415 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n352) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U418 ( .A(n353), .B(KEYINPUT89), .Z(n357) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n354), .B(G64GAT), .ZN(n435) );
  XNOR2_X1 U421 ( .A(n355), .B(n435), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n362) );
  XOR2_X1 U424 ( .A(G169GAT), .B(G8GAT), .Z(n420) );
  XNOR2_X1 U425 ( .A(n420), .B(n360), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n523) );
  XOR2_X1 U427 ( .A(n523), .B(KEYINPUT90), .Z(n363) );
  XNOR2_X1 U428 ( .A(n363), .B(KEYINPUT27), .ZN(n388) );
  XOR2_X1 U429 ( .A(n364), .B(KEYINPUT1), .Z(n366) );
  NAND2_X1 U430 ( .A1(G225GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n378) );
  XOR2_X1 U432 ( .A(KEYINPUT85), .B(KEYINPUT6), .Z(n368) );
  XNOR2_X1 U433 ( .A(G162GAT), .B(G85GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U435 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n370) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(KEYINPUT84), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U438 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U439 ( .A(G120GAT), .B(G148GAT), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n373), .B(G57GAT), .ZN(n436) );
  XNOR2_X1 U441 ( .A(n374), .B(n436), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n381) );
  INV_X1 U444 ( .A(n379), .ZN(n380) );
  XOR2_X1 U445 ( .A(n381), .B(n380), .Z(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT86), .B(n390), .ZN(n546) );
  INV_X1 U447 ( .A(n546), .ZN(n382) );
  AND2_X1 U448 ( .A1(n382), .A2(n530), .ZN(n383) );
  NAND2_X1 U449 ( .A1(n388), .A2(n383), .ZN(n533) );
  XNOR2_X1 U450 ( .A(n384), .B(KEYINPUT91), .ZN(n393) );
  NOR2_X1 U451 ( .A1(n534), .A2(n523), .ZN(n385) );
  NOR2_X1 U452 ( .A1(n472), .A2(n385), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n386), .B(KEYINPUT25), .ZN(n389) );
  NAND2_X1 U454 ( .A1(n472), .A2(n534), .ZN(n387) );
  XOR2_X1 U455 ( .A(n387), .B(KEYINPUT26), .Z(n574) );
  NAND2_X1 U456 ( .A1(n574), .A2(n388), .ZN(n545) );
  NAND2_X1 U457 ( .A1(n389), .A2(n545), .ZN(n391) );
  NAND2_X1 U458 ( .A1(n391), .A2(n390), .ZN(n392) );
  NAND2_X1 U459 ( .A1(n393), .A2(n392), .ZN(n395) );
  XOR2_X1 U460 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n397) );
  XNOR2_X1 U461 ( .A(G8GAT), .B(G64GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n413) );
  XOR2_X1 U463 ( .A(G57GAT), .B(G78GAT), .Z(n399) );
  XNOR2_X1 U464 ( .A(G155GAT), .B(G211GAT), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U466 ( .A(G71GAT), .B(KEYINPUT13), .Z(n434) );
  XOR2_X1 U467 ( .A(n400), .B(n434), .Z(n402) );
  XNOR2_X1 U468 ( .A(G183GAT), .B(G127GAT), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U470 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n404) );
  NAND2_X1 U471 ( .A1(G231GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U473 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U474 ( .A(G22GAT), .B(G15GAT), .Z(n408) );
  XNOR2_X1 U475 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U477 ( .A(G1GAT), .B(n409), .Z(n431) );
  XNOR2_X1 U478 ( .A(n431), .B(KEYINPUT14), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n413), .B(n412), .ZN(n562) );
  INV_X1 U481 ( .A(n562), .ZN(n586) );
  NOR2_X1 U482 ( .A1(n486), .A2(n586), .ZN(n414) );
  XOR2_X1 U483 ( .A(KEYINPUT96), .B(n414), .Z(n415) );
  NOR2_X1 U484 ( .A1(n590), .A2(n415), .ZN(n416) );
  XOR2_X1 U485 ( .A(KEYINPUT37), .B(n416), .Z(n518) );
  XOR2_X1 U486 ( .A(G197GAT), .B(G141GAT), .Z(n418) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G113GAT), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U489 ( .A(n419), .B(G50GAT), .Z(n422) );
  XNOR2_X1 U490 ( .A(n420), .B(G36GAT), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U492 ( .A(n423), .B(KEYINPUT29), .Z(n425) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U495 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U496 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n429) );
  XNOR2_X1 U497 ( .A(KEYINPUT68), .B(KEYINPUT70), .ZN(n428) );
  XNOR2_X1 U498 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U500 ( .A(n433), .B(n432), .Z(n579) );
  XOR2_X1 U501 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n441) );
  XNOR2_X1 U505 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U507 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U508 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n582) );
  NOR2_X1 U511 ( .A1(n480), .A2(n582), .ZN(n488) );
  NAND2_X1 U512 ( .A1(n518), .A2(n488), .ZN(n448) );
  NOR2_X1 U513 ( .A1(n530), .A2(n504), .ZN(n451) );
  INV_X1 U514 ( .A(G50GAT), .ZN(n449) );
  XOR2_X1 U515 ( .A(KEYINPUT41), .B(n582), .Z(n552) );
  INV_X1 U516 ( .A(n552), .ZN(n508) );
  INV_X1 U517 ( .A(n523), .ZN(n468) );
  INV_X1 U518 ( .A(KEYINPUT45), .ZN(n453) );
  XNOR2_X1 U519 ( .A(n453), .B(n452), .ZN(n454) );
  NOR2_X1 U520 ( .A1(n454), .A2(n582), .ZN(n455) );
  XOR2_X1 U521 ( .A(n455), .B(KEYINPUT108), .Z(n456) );
  NOR2_X1 U522 ( .A1(n579), .A2(n456), .ZN(n457) );
  XNOR2_X1 U523 ( .A(KEYINPUT109), .B(n457), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT47), .B(KEYINPUT107), .Z(n462) );
  NOR2_X1 U525 ( .A1(n480), .A2(n508), .ZN(n458) );
  XNOR2_X1 U526 ( .A(n458), .B(KEYINPUT46), .ZN(n459) );
  NOR2_X1 U527 ( .A1(n586), .A2(n459), .ZN(n460) );
  INV_X1 U528 ( .A(n559), .ZN(n568) );
  NAND2_X1 U529 ( .A1(n460), .A2(n568), .ZN(n461) );
  XOR2_X1 U530 ( .A(n462), .B(n461), .Z(n463) );
  AND2_X1 U531 ( .A1(n464), .A2(n463), .ZN(n467) );
  NAND2_X1 U532 ( .A1(n468), .A2(n548), .ZN(n470) );
  XOR2_X1 U533 ( .A(KEYINPUT116), .B(KEYINPUT54), .Z(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U535 ( .A1(n546), .A2(n471), .ZN(n576) );
  NOR2_X1 U536 ( .A1(n472), .A2(n576), .ZN(n474) );
  XNOR2_X1 U537 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n474), .B(n473), .ZN(n476) );
  NAND2_X1 U539 ( .A1(n476), .A2(n475), .ZN(n567) );
  NOR2_X1 U540 ( .A1(n508), .A2(n567), .ZN(n479) );
  XNOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n477) );
  INV_X1 U542 ( .A(G169GAT), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT118), .B(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1348GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n485) );
  NAND2_X1 U546 ( .A1(n586), .A2(n568), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(n487) );
  NOR2_X1 U548 ( .A1(n487), .A2(n486), .ZN(n509) );
  NAND2_X1 U549 ( .A1(n509), .A2(n488), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT93), .B(n489), .Z(n496) );
  NOR2_X1 U551 ( .A1(n546), .A2(n496), .ZN(n490) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(n490), .Z(n491) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U554 ( .A1(n523), .A2(n496), .ZN(n492) );
  XOR2_X1 U555 ( .A(G8GAT), .B(n492), .Z(G1325GAT) );
  NOR2_X1 U556 ( .A1(n534), .A2(n496), .ZN(n494) );
  XNOR2_X1 U557 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  NOR2_X1 U560 ( .A1(n530), .A2(n496), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(KEYINPUT95), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(G1327GAT) );
  NOR2_X1 U563 ( .A1(n504), .A2(n546), .ZN(n501) );
  XOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U565 ( .A(KEYINPUT97), .B(n499), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n504), .A2(n523), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT98), .B(n502), .Z(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT99), .ZN(n506) );
  NOR2_X1 U571 ( .A1(n534), .A2(n504), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U574 ( .A1(n508), .A2(n579), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n519), .A2(n509), .ZN(n515) );
  NOR2_X1 U576 ( .A1(n546), .A2(n515), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(KEYINPUT101), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n523), .A2(n515), .ZN(n513) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n534), .A2(n515), .ZN(n514) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n530), .A2(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U588 ( .A1(n546), .A2(n529), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n521), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(KEYINPUT103), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT104), .B(n524), .Z(n525) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n534), .A2(n529), .ZN(n526) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n528) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(KEYINPUT106), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n532) );
  NOR2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(n532), .B(n531), .Z(G1339GAT) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n548), .A2(n535), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT111), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n579), .A2(n542), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U606 ( .A1(n542), .A2(n552), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n542), .A2(n586), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U612 ( .A1(n542), .A2(n559), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT113), .Z(n551) );
  NOR2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT112), .B(n549), .Z(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n579), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT114), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U622 ( .A1(n560), .A2(n552), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT115), .Z(n558) );
  NAND2_X1 U626 ( .A1(n586), .A2(n560), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n562), .A2(n567), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT119), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT120), .B(KEYINPUT58), .Z(n566) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n566), .B(n565), .ZN(n570) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(n570), .B(n569), .Z(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n572) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT123), .B(n573), .Z(n581) );
  INV_X1 U642 ( .A(n574), .ZN(n575) );
  NOR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n578) );
  INV_X1 U644 ( .A(KEYINPUT122), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n587), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n584) );
  NAND2_X1 U649 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT126), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

