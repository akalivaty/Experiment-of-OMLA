//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G143), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI211_X1 g007(.A(G128), .B(new_n191), .C1(new_n192), .C2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n195), .B1(new_n192), .B2(new_n193), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n198));
  OAI22_X1  g012(.A1(new_n194), .A2(KEYINPUT1), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(new_n193), .ZN(new_n205));
  INV_X1    g019(.A(new_n195), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n208), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n202), .A2(new_n204), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n190), .B1(new_n214), .B2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n209), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n201), .B1(new_n218), .B2(new_n200), .ZN(new_n219));
  INV_X1    g033(.A(G224), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G953), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n219), .B(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(G110), .B(G122), .Z(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT80), .B(G104), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT80), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G104), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n231), .A3(new_n226), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n228), .A2(KEYINPUT3), .A3(G107), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(G104), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n228), .A2(KEYINPUT80), .ZN(new_n237));
  OAI211_X1 g051(.A(KEYINPUT81), .B(G107), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n227), .A2(new_n233), .A3(new_n235), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n227), .A4(new_n238), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n245));
  INV_X1    g059(.A(G113), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT2), .A3(G113), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n247), .A2(new_n249), .B1(new_n245), .B2(new_n246), .ZN(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G119), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n250), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n239), .A2(new_n256), .A3(G101), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n244), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT85), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n232), .B1(G104), .B2(new_n226), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G101), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n243), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n265));
  INV_X1    g079(.A(G119), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G116), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(G113), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT84), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n250), .A2(new_n251), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n258), .A2(new_n259), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n259), .B1(new_n258), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n223), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n223), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n258), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT6), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT6), .B(new_n223), .C1(new_n272), .C2(new_n273), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n222), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n219), .B(KEYINPUT7), .C1(new_n220), .C2(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n262), .A3(new_n270), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n223), .B(KEYINPUT8), .Z(new_n283));
  AND2_X1   g097(.A1(new_n270), .A2(new_n268), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n282), .B(new_n283), .C1(new_n262), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n286));
  OAI221_X1 g100(.A(new_n201), .B1(new_n286), .B2(new_n221), .C1(new_n218), .C2(new_n200), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n281), .A2(new_n276), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n188), .B1(new_n280), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n258), .A2(new_n271), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT85), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n258), .A2(new_n271), .A3(new_n259), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n275), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n277), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n279), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n222), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n290), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n187), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n291), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(G952), .ZN(new_n305));
  AOI211_X1 g119(.A(G953), .B(new_n305), .C1(G234), .C2(G237), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT73), .B(G902), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n308), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT21), .B(G898), .Z(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT95), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n307), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n299), .A2(KEYINPUT86), .A3(new_n187), .A4(new_n300), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n303), .A2(new_n304), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n308), .A3(G143), .A4(G214), .ZN(new_n319));
  INV_X1    g133(.A(G214), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(G237), .A3(G953), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT87), .B(new_n319), .C1(new_n192), .C2(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n319), .A2(KEYINPUT87), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(G131), .A3(new_n323), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n200), .A2(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT16), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n336), .A2(new_n331), .A3(KEYINPUT77), .A4(G125), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n193), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n333), .A2(new_n335), .A3(G146), .A4(new_n337), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n322), .A2(G131), .A3(new_n323), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n329), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n324), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n322), .A2(KEYINPUT18), .A3(G131), .A4(new_n323), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n332), .A2(new_n334), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(new_n193), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n326), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G113), .B(G122), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(new_n228), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n345), .A2(new_n354), .A3(new_n351), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n289), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G475), .ZN(new_n360));
  AND2_X1   g174(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n332), .B(new_n334), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(new_n193), .C1(new_n349), .C2(new_n362), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n364), .A2(new_n340), .ZN(new_n365));
  AOI21_X1  g179(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n343), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n351), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n355), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(KEYINPUT89), .A3(new_n355), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n357), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n374));
  NOR2_X1   g188(.A1(G475), .A2(G902), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n373), .A2(KEYINPUT90), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n360), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n357), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT89), .B1(new_n368), .B2(new_n355), .ZN(new_n379));
  AOI211_X1 g193(.A(new_n370), .B(new_n354), .C1(new_n351), .C2(new_n367), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n375), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT20), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT9), .B(G234), .Z(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(new_n391), .A3(G953), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT13), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n192), .B2(new_n197), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT91), .B1(new_n189), .B2(G128), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n197), .A3(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n203), .A2(G143), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT13), .B(G128), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT92), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(G134), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n403), .B2(G134), .ZN(new_n406));
  XNOR2_X1  g220(.A(G116), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n226), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n214), .A2(G128), .ZN(new_n409));
  OR2_X1    g223(.A1(KEYINPUT66), .A2(G134), .ZN(new_n410));
  NAND2_X1  g224(.A1(KEYINPUT66), .A2(G134), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n412), .A3(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n405), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n399), .ZN(new_n416));
  AND2_X1   g230(.A1(KEYINPUT66), .A2(G134), .ZN(new_n417));
  NOR2_X1   g231(.A1(KEYINPUT66), .A2(G134), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n407), .A2(new_n226), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n407), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G122), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n425), .A2(G116), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n424), .B(G107), .C1(new_n423), .C2(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n421), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n393), .B1(new_n415), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n403), .A2(G134), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT92), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n403), .A2(new_n404), .A3(G134), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n413), .A3(new_n408), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n421), .A2(new_n422), .A3(new_n427), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n392), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(KEYINPUT93), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n433), .A2(new_n437), .A3(new_n434), .A4(new_n392), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n310), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G478), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n436), .A2(new_n310), .A3(new_n438), .A4(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n388), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G469), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT1), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n215), .A2(new_n452), .A3(G128), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n215), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n192), .B2(new_n193), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n197), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n215), .A2(KEYINPUT82), .A3(new_n452), .A4(G128), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n263), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n410), .A2(G137), .A3(new_n411), .ZN(new_n465));
  NOR2_X1   g279(.A1(G134), .A2(G137), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n464), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NOR4_X1   g282(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT11), .A4(G137), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n325), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G137), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n419), .A2(new_n464), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n466), .B1(new_n419), .B2(G137), .ZN(new_n473));
  OAI211_X1 g287(.A(G131), .B(new_n472), .C1(new_n473), .C2(new_n464), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n210), .A2(new_n211), .B1(new_n216), .B2(new_n215), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n244), .A2(new_n213), .A3(new_n476), .A4(new_n257), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n263), .A2(KEYINPUT10), .A3(new_n199), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n463), .A2(new_n475), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n262), .B(new_n453), .C1(new_n196), .C2(new_n198), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n461), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n470), .A2(new_n474), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n482), .A2(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT12), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G140), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n308), .A2(G227), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n488), .B(new_n489), .Z(new_n490));
  AND4_X1   g304(.A1(new_n479), .A2(new_n485), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n463), .A2(new_n477), .A3(new_n478), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n482), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n490), .B1(new_n493), .B2(new_n479), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n451), .B(new_n310), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(G469), .A2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n479), .A3(new_n487), .ZN(new_n497));
  INV_X1    g311(.A(new_n490), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n479), .A3(new_n490), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(G469), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n317), .A2(new_n450), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n266), .A2(G128), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n197), .A2(G119), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(KEYINPUT76), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G110), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n511));
  OAI211_X1 g325(.A(G119), .B(new_n197), .C1(new_n511), .C2(KEYINPUT23), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n506), .B(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n515), .A2(new_n508), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT24), .B(G110), .Z(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT78), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n349), .A2(new_n193), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n340), .A4(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n513), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n517), .B1(new_n515), .B2(new_n508), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n340), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT78), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n516), .A2(new_n517), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n509), .A2(new_n512), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n526), .B(new_n341), .C1(new_n510), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT22), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(G137), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n521), .A2(new_n525), .A3(new_n528), .A4(new_n532), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT25), .B1(new_n536), .B2(new_n309), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n391), .B1(new_n310), .B2(G234), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n534), .A2(new_n539), .A3(new_n310), .A4(new_n535), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n538), .A2(G902), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n534), .A2(new_n542), .A3(new_n535), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n482), .A2(new_n476), .A3(new_n213), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT67), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n471), .A2(G134), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n419), .B2(new_n471), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n549), .B2(new_n325), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n412), .A2(G137), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT67), .B(G131), .C1(new_n551), .C2(new_n548), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n199), .A2(new_n470), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n545), .A2(new_n546), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n546), .B1(new_n545), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n255), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n545), .A2(new_n254), .A3(new_n553), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n318), .A2(new_n308), .A3(G210), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT71), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT72), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT31), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n565), .B2(KEYINPUT31), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n553), .B1(new_n475), .B2(new_n218), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n255), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n569), .B1(new_n571), .B2(new_n557), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n557), .A2(new_n569), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n563), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n556), .A2(new_n576), .A3(new_n557), .A4(new_n564), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n567), .A2(new_n568), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(G472), .A2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT32), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n565), .A2(KEYINPUT31), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT72), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n575), .A2(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT31), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n580), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n545), .A2(new_n254), .A3(new_n553), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n254), .B1(new_n545), .B2(new_n553), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT28), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n573), .A3(new_n564), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n570), .A2(KEYINPUT30), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n545), .A2(new_n546), .A3(new_n553), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n591), .B1(new_n598), .B2(new_n255), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n594), .B(new_n595), .C1(new_n599), .C2(new_n564), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n593), .A2(KEYINPUT29), .A3(new_n573), .A4(new_n564), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n310), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT74), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(KEYINPUT74), .A3(G472), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT79), .B(new_n544), .C1(new_n590), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT79), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n579), .A2(KEYINPUT32), .A3(new_n581), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n588), .B1(new_n587), .B2(new_n580), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n602), .A2(KEYINPUT74), .A3(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT74), .B1(new_n602), .B2(G472), .ZN(new_n613));
  OAI22_X1  g427(.A1(new_n610), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n544), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n505), .B1(new_n608), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(new_n504), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n579), .B2(new_n309), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n587), .A2(new_n580), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n615), .A4(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n187), .B1(new_n299), .B2(new_n300), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n188), .B(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n304), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n315), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n439), .A2(new_n440), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n436), .A2(new_n629), .A3(new_n438), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n429), .A2(KEYINPUT33), .A3(new_n435), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n310), .A2(G478), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n387), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n626), .A2(new_n627), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n623), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(G475), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n358), .B2(new_n289), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n383), .B2(new_n385), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n446), .A2(new_n448), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n626), .A2(new_n627), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n623), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n620), .A2(new_n621), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n529), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n542), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n541), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n650), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n655), .B(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(KEYINPUT98), .A3(new_n621), .A4(new_n620), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n505), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT37), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n510), .ZN(G12));
  AOI21_X1  g477(.A(new_n656), .B1(new_n590), .B2(new_n607), .ZN(new_n664));
  INV_X1    g478(.A(new_n304), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n291), .B2(new_n301), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n307), .B1(new_n312), .B2(G900), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT99), .Z(new_n668));
  NOR2_X1   g482(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT100), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n666), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n664), .A2(new_n619), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NOR2_X1   g489(.A1(new_n599), .A2(new_n563), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n591), .A2(new_n592), .ZN(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n677), .B2(new_n563), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n590), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n668), .B(KEYINPUT39), .Z(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n504), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n665), .B(new_n682), .C1(KEYINPUT40), .C2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n303), .A2(new_n316), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT38), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n387), .A2(new_n644), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n687), .A2(new_n541), .A3(new_n692), .A4(new_n654), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n192), .ZN(G45));
  INV_X1    g508(.A(new_n668), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n387), .A2(new_n634), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n664), .A2(new_n619), .A3(new_n666), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  OAI21_X1  g512(.A(new_n310), .B1(new_n491), .B2(new_n494), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n503), .A3(new_n495), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n636), .A2(new_n614), .A3(new_n615), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n544), .B1(new_n590), .B2(new_n607), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n636), .A4(new_n702), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT41), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G113), .ZN(G15));
  NAND4_X1  g524(.A1(new_n646), .A2(new_n614), .A3(new_n615), .A4(new_n702), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT102), .B(G116), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G18));
  NOR2_X1   g527(.A1(new_n450), .A2(new_n627), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n626), .A2(new_n701), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n614), .A2(new_n714), .A3(new_n715), .A4(new_n659), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  AOI21_X1  g531(.A(new_n576), .B1(new_n599), .B2(new_n564), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n580), .B1(new_n578), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(KEYINPUT103), .B(new_n580), .C1(new_n578), .C2(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(G472), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n587), .B2(new_n310), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n723), .A2(new_n725), .A3(new_n544), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n701), .A2(new_n627), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n691), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n387), .A2(KEYINPUT104), .A3(new_n644), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n666), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n626), .B1(new_n730), .B2(new_n731), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n726), .A3(new_n736), .A4(new_n727), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  AND2_X1   g553(.A1(new_n721), .A2(new_n722), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n696), .A3(new_n620), .A4(new_n655), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n702), .A2(new_n666), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n200), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n610), .B2(new_n611), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n582), .A2(KEYINPUT108), .A3(new_n589), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n607), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n496), .B(KEYINPUT106), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n495), .A2(new_n501), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n503), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n665), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND4_X1   g568(.A1(KEYINPUT42), .A2(new_n387), .A3(new_n634), .A4(new_n695), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n688), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n748), .A2(new_n756), .A3(new_n615), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n748), .A2(new_n756), .A3(KEYINPUT109), .A4(new_n615), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n753), .B1(new_n316), .B2(new_n303), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n705), .A2(new_n696), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n759), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n614), .A3(new_n615), .A4(new_n669), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  AOI21_X1  g582(.A(new_n665), .B1(new_n303), .B2(new_n316), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n388), .A2(new_n634), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT43), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n651), .A3(new_n655), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n499), .A2(new_n500), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT45), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(G469), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n749), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT110), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  INV_X1    g595(.A(new_n495), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n783), .A2(KEYINPUT111), .A3(new_n751), .A4(new_n684), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n779), .A2(new_n780), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n781), .A2(new_n782), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n751), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n785), .B1(new_n788), .B2(new_n683), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n769), .B(new_n773), .C1(new_n784), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  AOI22_X1  g605(.A1(new_n582), .A2(new_n589), .B1(new_n605), .B2(new_n606), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n696), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n783), .B2(new_n751), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n544), .A3(new_n769), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  AND3_X1   g613(.A1(new_n759), .A2(new_n760), .A3(new_n764), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n711), .A2(new_n716), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n723), .A2(new_n725), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n761), .A2(new_n655), .A3(new_n696), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n767), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n708), .A2(new_n738), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n388), .A2(new_n644), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n622), .A2(new_n317), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n303), .A2(new_n315), .A3(new_n316), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n810));
  INV_X1    g624(.A(new_n635), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n304), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT113), .B1(new_n317), .B2(new_n635), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n623), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n617), .A2(new_n661), .A3(new_n808), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n643), .A2(new_n449), .A3(new_n695), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n643), .A2(new_n449), .A3(new_n818), .A4(new_n695), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n820), .A2(new_n769), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n820), .B2(new_n769), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n504), .B(new_n656), .C1(new_n590), .C2(new_n607), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n688), .A2(new_n304), .A3(new_n817), .A4(new_n819), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n820), .A2(new_n769), .A3(new_n821), .ZN(new_n831));
  AND4_X1   g645(.A1(KEYINPUT116), .A2(new_n825), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n815), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n806), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n711), .A2(new_n716), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n737), .B2(new_n734), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n765), .A2(new_n838), .A3(new_n708), .A4(new_n804), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n622), .A2(new_n317), .A3(new_n807), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n705), .A2(new_n609), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT79), .B1(new_n792), .B2(new_n544), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n843), .B2(new_n505), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n814), .A2(new_n661), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT116), .B1(new_n824), .B2(new_n825), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n832), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n741), .A2(new_n742), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n668), .A2(new_n751), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n750), .A2(new_n541), .A3(new_n654), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n735), .A2(new_n681), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n674), .A2(new_n697), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n671), .A2(new_n673), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n743), .B1(new_n857), .B2(new_n825), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(KEYINPUT52), .A3(new_n697), .A4(new_n853), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT119), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n849), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n697), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n853), .A2(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n674), .A2(new_n850), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n856), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n806), .A2(new_n834), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n305), .A2(G953), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n700), .A2(new_n495), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n751), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n795), .A2(new_n796), .A3(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n771), .A2(new_n306), .A3(new_n726), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(new_n769), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n769), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n544), .A3(new_n701), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n306), .A3(new_n682), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n889), .A2(new_n387), .A3(new_n634), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n884), .A2(new_n665), .A3(new_n689), .A4(new_n702), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT50), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n306), .A2(new_n771), .A3(new_n702), .A4(new_n769), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n802), .A2(new_n655), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n886), .A2(new_n890), .A3(new_n893), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n748), .A2(new_n615), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT48), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n883), .A2(new_n885), .B1(new_n895), .B2(new_n894), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT51), .A3(new_n890), .A4(new_n893), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n880), .A2(new_n899), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n849), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n872), .B2(new_n873), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n861), .A2(new_n863), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n848), .B2(new_n836), .ZN(new_n910));
  OAI221_X1 g724(.A(KEYINPUT54), .B1(new_n906), .B2(new_n908), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n889), .A2(new_n635), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n879), .A2(new_n905), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n884), .A2(new_n715), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT120), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n913), .A2(new_n915), .B1(G952), .B2(G953), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT49), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n615), .B1(new_n881), .B2(new_n917), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n918), .A2(new_n751), .A3(new_n665), .A4(new_n770), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n881), .A2(new_n917), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n682), .A3(new_n689), .A4(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT112), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n916), .A2(new_n922), .ZN(G75));
  OAI22_X1  g737(.A1(new_n910), .A2(KEYINPUT53), .B1(new_n875), .B2(new_n874), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n309), .A3(new_n188), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT121), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n297), .B(new_n298), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n929), .ZN(new_n931));
  AOI211_X1 g745(.A(KEYINPUT121), .B(new_n931), .C1(new_n925), .C2(new_n926), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n925), .A2(KEYINPUT121), .A3(new_n926), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n305), .A2(G953), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT122), .Z(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT123), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n930), .A2(new_n932), .A3(new_n937), .ZN(G51));
  INV_X1    g752(.A(new_n935), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n749), .A2(KEYINPUT57), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n749), .A2(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n877), .A2(new_n878), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n924), .A2(KEYINPUT54), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n491), .A2(new_n494), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n924), .A2(G469), .A3(new_n309), .A4(new_n775), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n939), .B1(new_n946), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n309), .B(new_n949), .C1(new_n865), .C2(new_n876), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n373), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n924), .A2(new_n309), .A3(new_n381), .A4(new_n949), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n935), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n935), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G60));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n879), .B2(new_n911), .ZN(new_n961));
  INV_X1    g775(.A(new_n632), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n936), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n942), .B2(new_n943), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n960), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT125), .Z(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT60), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n536), .B1(new_n877), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n924), .A2(new_n653), .A3(new_n969), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n936), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G66));
  AOI21_X1  g789(.A(new_n308), .B1(new_n314), .B2(G224), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n838), .A2(new_n845), .A3(new_n844), .A4(new_n708), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(new_n308), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n278), .B(new_n279), .C1(G898), .C2(new_n308), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT127), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  OAI21_X1  g796(.A(new_n363), .B1(new_n349), .B2(new_n362), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n598), .B(new_n983), .Z(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n798), .A2(new_n790), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n866), .B1(new_n868), .B2(new_n871), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n765), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n735), .B(new_n900), .C1(new_n784), .C2(new_n789), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n986), .A2(new_n767), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n984), .B(new_n985), .C1(new_n990), .C2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n693), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT62), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n887), .B1(new_n635), .B2(new_n807), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n843), .A2(new_n685), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n986), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n997), .A2(new_n308), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n991), .B1(new_n998), .B2(new_n984), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n308), .B1(G227), .B2(G900), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n997), .B2(new_n978), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n939), .B1(new_n1004), .B2(new_n676), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n990), .B2(new_n978), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n563), .A3(new_n599), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n599), .B(new_n564), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1009));
  OAI221_X1 g823(.A(new_n1009), .B1(new_n906), .B2(new_n908), .C1(new_n907), .C2(new_n910), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1005), .A2(new_n1007), .A3(new_n1010), .ZN(G57));
endmodule


