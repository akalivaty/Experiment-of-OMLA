//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(G85gat), .ZN(new_n202));
  INV_X1    g001(.A(G92gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT90), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G99gat), .B(G106gat), .Z(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(KEYINPUT92), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(KEYINPUT91), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(KEYINPUT91), .B2(new_n212), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n206), .A2(KEYINPUT90), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n205), .A3(new_n207), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n209), .A2(KEYINPUT92), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n222), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT14), .B(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G43gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n227), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n231), .B2(new_n232), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT93), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n221), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n234), .B2(new_n236), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n238), .B(new_n239), .C1(new_n241), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n247));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n239), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n221), .B(KEYINPUT93), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n248), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT95), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n255), .A3(KEYINPUT94), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G134gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(G162gat), .Z(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n257), .B1(new_n258), .B2(new_n261), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G57gat), .B(G64gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G78gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G127gat), .B(G155gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT89), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n275), .B(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G183gat), .B(G211gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G15gat), .B(G22gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT16), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(G1gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(G1gat), .B2(new_n281), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(G8gat), .Z(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n272), .B2(new_n271), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n280), .B(new_n288), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n221), .A2(new_n270), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT10), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n219), .A2(new_n220), .A3(new_n271), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n270), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n297), .B(KEYINPUT96), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n291), .B2(new_n293), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT97), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G120gat), .B(G148gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G176gat), .B(G204gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n301), .B2(new_n302), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n300), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n298), .B1(new_n294), .B2(new_n295), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n310), .B2(new_n301), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(G197gat), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT11), .B(G169gat), .Z(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n316), .B(KEYINPUT12), .Z(new_n317));
  INV_X1    g116(.A(new_n285), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(new_n237), .ZN(new_n319));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT13), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n242), .B2(new_n244), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n237), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n320), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n322), .B1(new_n327), .B2(KEYINPUT18), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n320), .B(new_n324), .C1(new_n245), .C2(new_n318), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT18), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n317), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n335));
  INV_X1    g134(.A(new_n317), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(new_n322), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(KEYINPUT88), .B(new_n317), .C1(new_n328), .C2(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n290), .A2(new_n312), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G15gat), .B(G43gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G127gat), .ZN(new_n349));
  INV_X1    g148(.A(G127gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G134gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT70), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G113gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G120gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n349), .B2(new_n351), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n357), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n350), .A2(G134gat), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n366), .A2(new_n363), .B1(KEYINPUT68), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n351), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n360), .A2(new_n365), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G169gat), .ZN(new_n376));
  INV_X1    g175(.A(G176gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT23), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(G169gat), .B2(G176gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT27), .B(G183gat), .ZN(new_n384));
  INV_X1    g183(.A(G190gat), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT28), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G183gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT27), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G183gat), .ZN(new_n390));
  AND4_X1   g189(.A1(KEYINPUT28), .A2(new_n388), .A3(new_n390), .A4(new_n385), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OR3_X1    g194(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n383), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT67), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(G183gat), .B2(G190gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n398), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT66), .ZN(new_n408));
  INV_X1    g207(.A(new_n372), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n373), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n405), .A2(new_n408), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n378), .B(new_n380), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n401), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n371), .B1(new_n400), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT64), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n412), .A2(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT25), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n375), .A2(new_n382), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n388), .A2(new_n390), .A3(new_n385), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT28), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n384), .A2(KEYINPUT28), .A3(new_n385), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n395), .A2(new_n396), .B1(G183gat), .B2(G190gat), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n367), .A2(KEYINPUT68), .ZN(new_n431));
  XNOR2_X1  g230(.A(G113gat), .B(G120gat), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n370), .B(new_n431), .C1(KEYINPUT1), .C2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n362), .B(new_n363), .C1(new_n434), .C2(new_n352), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n353), .A2(new_n359), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n420), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n347), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n420), .B1(new_n418), .B2(new_n438), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT34), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI211_X1 g243(.A(KEYINPUT34), .B(new_n420), .C1(new_n418), .C2(new_n438), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n449));
  INV_X1    g248(.A(new_n439), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n447), .A2(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n444), .A2(new_n445), .ZN(new_n452));
  INV_X1    g251(.A(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n450), .A2(new_n449), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n446), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n451), .A2(KEYINPUT36), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT36), .B1(new_n451), .B2(new_n456), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(G57gat), .B(G85gat), .Z(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT78), .ZN(new_n461));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n463), .B(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n467));
  NAND2_X1  g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT2), .ZN(new_n469));
  OR2_X1    g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(G141gat), .A2(G148gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G155gat), .B(G162gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(KEYINPUT74), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n472), .B2(new_n474), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G141gat), .B(G148gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT2), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(G155gat), .B2(G162gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n473), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT3), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n477), .A2(new_n485), .A3(new_n437), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT76), .A4(new_n437), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G225gat), .A2(G233gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n475), .A2(new_n476), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n437), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n483), .A2(new_n484), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n491), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n371), .A2(new_n495), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n493), .A2(new_n437), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n497), .B1(new_n488), .B2(new_n489), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n491), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n466), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(new_n466), .A3(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT79), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n511), .B(new_n512), .C1(new_n509), .C2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n463), .B(new_n464), .ZN(new_n515));
  AND4_X1   g314(.A1(new_n507), .A2(new_n490), .A3(new_n491), .A4(new_n498), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n506), .B2(new_n491), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT79), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n510), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G8gat), .B(G36gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n522), .B(new_n523), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n400), .B2(new_n417), .ZN(new_n528));
  NAND2_X1  g327(.A1(G211gat), .A2(G218gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT22), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(G197gat), .A2(G204gat), .ZN(new_n532));
  AND2_X1   g331(.A1(G197gat), .A2(G204gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(G211gat), .A2(G218gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n529), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n534), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G226gat), .A2(G233gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n422), .A2(new_n430), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n528), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(new_n528), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n525), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n422), .A2(new_n430), .A3(new_n540), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n526), .B1(new_n422), .B2(new_n430), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n539), .A3(new_n541), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n524), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(KEYINPUT30), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n547), .A2(new_n551), .A3(new_n548), .A4(new_n524), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n521), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n467), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n483), .B2(new_n484), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n538), .B1(new_n557), .B2(KEYINPUT29), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n535), .A2(new_n529), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT29), .B1(new_n534), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n532), .ZN(new_n561));
  NAND2_X1  g360(.A1(G197gat), .A2(G204gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n561), .A2(new_n562), .B1(new_n530), .B2(new_n529), .ZN(new_n563));
  INV_X1    g362(.A(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(KEYINPUT81), .B(new_n493), .C1(new_n566), .C2(new_n556), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT81), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n556), .B1(new_n560), .B2(new_n565), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(new_n495), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n558), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G228gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT3), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n538), .B2(KEYINPUT29), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n573), .B1(new_n576), .B2(new_n493), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n558), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G22gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n571), .A2(new_n573), .B1(new_n577), .B2(new_n558), .ZN(new_n581));
  INV_X1    g380(.A(G22gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G78gat), .B(G106gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G50gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT80), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n581), .A2(KEYINPUT83), .A3(new_n582), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT83), .B1(new_n581), .B2(new_n582), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n579), .A2(KEYINPUT82), .A3(G22gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT82), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n581), .B2(new_n582), .ZN(new_n595));
  INV_X1    g394(.A(new_n587), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n589), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n459), .B1(new_n555), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n519), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n509), .A2(KEYINPUT84), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n553), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n491), .B1(new_n490), .B2(new_n498), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n515), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n501), .A2(new_n502), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n609), .B2(new_n491), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n506), .B2(new_n491), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n608), .B1(new_n607), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT85), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n512), .A2(new_n511), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n602), .A3(new_n603), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n547), .A2(new_n548), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n525), .B1(new_n618), .B2(KEYINPUT37), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n547), .B2(new_n548), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT38), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n525), .A2(KEYINPUT37), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n544), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n620), .B1(new_n543), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n547), .A2(KEYINPUT86), .A3(new_n548), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n622), .A2(new_n630), .A3(new_n549), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n617), .A2(new_n510), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n505), .A2(new_n508), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT84), .B1(new_n633), .B2(new_n515), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n601), .B(new_n466), .C1(new_n505), .C2(new_n508), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT85), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n605), .A2(new_n606), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n466), .A3(new_n611), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n636), .A2(new_n637), .A3(new_n642), .A4(new_n553), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n615), .A2(new_n632), .A3(new_n643), .A4(new_n598), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n598), .A2(new_n554), .A3(new_n456), .A4(new_n451), .ZN(new_n645));
  INV_X1    g444(.A(new_n510), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n513), .B1(new_n633), .B2(new_n515), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n512), .A2(new_n511), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n509), .A2(new_n513), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT35), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  AND4_X1   g451(.A1(new_n598), .A2(new_n554), .A3(new_n456), .A4(new_n451), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT35), .B1(new_n617), .B2(new_n510), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n600), .A2(new_n644), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n341), .A2(KEYINPUT98), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT98), .B1(new_n341), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n651), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g462(.A(G8gat), .B1(new_n660), .B2(new_n554), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n660), .A2(new_n554), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n668), .A2(KEYINPUT99), .A3(new_n665), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT99), .B1(new_n668), .B2(new_n665), .ZN(new_n670));
  OAI221_X1 g469(.A(new_n664), .B1(new_n665), .B2(new_n668), .C1(new_n669), .C2(new_n670), .ZN(G1325gat));
  INV_X1    g470(.A(new_n459), .ZN(new_n672));
  OAI21_X1  g471(.A(G15gat), .B1(new_n660), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n454), .A2(new_n455), .A3(new_n446), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n455), .B1(new_n454), .B2(new_n446), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G15gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n673), .B1(new_n660), .B2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n660), .A2(new_n598), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n555), .A2(new_n599), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n644), .A2(new_n684), .A3(new_n672), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n652), .A2(new_n655), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n265), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(KEYINPUT100), .B(KEYINPUT44), .C1(new_n656), .C2(new_n265), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n264), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n262), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n685), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n600), .A2(KEYINPUT101), .A3(new_n644), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n652), .A2(new_n655), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n652), .B2(new_n655), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n688), .B(new_n693), .C1(new_n697), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n289), .A2(new_n340), .A3(new_n312), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n521), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n687), .A2(new_n704), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n222), .A3(new_n651), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(G1328gat));
  OAI21_X1  g509(.A(G36gat), .B1(new_n705), .B2(new_n554), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n712));
  AOI21_X1  g511(.A(G36gat), .B1(new_n712), .B2(KEYINPUT46), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n707), .A2(new_n553), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  OAI21_X1  g517(.A(G43gat), .B1(new_n705), .B2(new_n672), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n707), .A2(new_n721), .A3(new_n676), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n722), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n719), .A2(KEYINPUT105), .A3(KEYINPUT47), .A4(new_n722), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(new_n730), .ZN(G1330gat));
  NOR3_X1   g530(.A1(new_n705), .A2(new_n229), .A3(new_n598), .ZN(new_n732));
  AOI21_X1  g531(.A(G50gat), .B1(new_n707), .B2(new_n599), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT48), .Z(G1331gat));
  OAI211_X1 g534(.A(new_n695), .B(new_n696), .C1(new_n700), .C2(new_n699), .ZN(new_n736));
  INV_X1    g535(.A(new_n340), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n290), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n736), .A2(new_n312), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n651), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g540(.A(new_n739), .B(KEYINPUT106), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n553), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n743), .B2(new_n744), .ZN(G1333gat));
  AOI21_X1  g546(.A(G71gat), .B1(new_n739), .B2(new_n676), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n459), .A2(G71gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n742), .A2(new_n599), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n289), .A2(new_n737), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n312), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT108), .B1(new_n703), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n760), .B(new_n756), .C1(new_n691), .C2(new_n702), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n521), .ZN(new_n764));
  INV_X1    g563(.A(new_n312), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n693), .B(new_n755), .C1(new_n697), .C2(new_n701), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n693), .A4(new_n755), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n202), .A3(new_n651), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n764), .A2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n768), .A2(new_n773), .A3(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n766), .A2(KEYINPUT109), .A3(new_n767), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n554), .A2(G92gat), .ZN(new_n776));
  AND4_X1   g575(.A1(new_n312), .A2(new_n774), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n762), .A3(new_n553), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(G92gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n756), .B1(new_n691), .B2(new_n702), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n553), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n781), .B1(new_n783), .B2(G92gat), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n776), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n779), .A2(new_n780), .B1(new_n787), .B2(new_n788), .ZN(G1337gat));
  XNOR2_X1  g588(.A(KEYINPUT112), .B(G99gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n676), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n763), .A2(new_n672), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n790), .ZN(G1338gat));
  INV_X1    g592(.A(G106gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n599), .A2(new_n794), .A3(new_n312), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n774), .A2(KEYINPUT113), .A3(new_n775), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n774), .A2(new_n775), .A3(new_n796), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n758), .A2(new_n761), .A3(new_n598), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n797), .B(new_n800), .C1(new_n801), .C2(new_n794), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n794), .B1(new_n782), .B2(new_n599), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n795), .B1(new_n768), .B2(new_n769), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1339gat));
  INV_X1    g606(.A(new_n289), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n294), .A2(new_n298), .A3(new_n295), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n300), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n306), .B1(new_n310), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n309), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n812), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n813), .A2(KEYINPUT114), .A3(new_n309), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n339), .A3(new_n338), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n326), .B1(new_n323), .B2(new_n325), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n319), .B2(new_n321), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n316), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n312), .A2(new_n337), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n693), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n337), .A2(new_n823), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n263), .B2(new_n264), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n818), .A2(new_n819), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n808), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n738), .A2(new_n765), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n521), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n653), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n737), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n312), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n289), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g640(.A1(new_n676), .A2(new_n598), .ZN(new_n842));
  NOR4_X1   g641(.A1(new_n265), .A2(G134gat), .A3(new_n553), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n834), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT56), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n348), .B1(new_n835), .B2(new_n693), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  NOR2_X1   g646(.A1(new_n459), .A2(new_n521), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n554), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT116), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n693), .A2(new_n819), .A3(new_n818), .A4(new_n828), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n817), .A2(new_n816), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n309), .A3(new_n813), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n824), .B1(new_n340), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n265), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n289), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n290), .A2(new_n312), .A3(new_n737), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n599), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n850), .B1(new_n858), .B2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n832), .A2(new_n833), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n599), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n737), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G141gat), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n598), .B1(new_n832), .B2(new_n833), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n848), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n553), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n340), .A2(G141gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n864), .B2(new_n869), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n863), .B2(G141gat), .ZN(new_n873));
  OAI22_X1  g672(.A1(new_n871), .A2(new_n872), .B1(KEYINPUT58), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n864), .A2(new_n869), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n874), .A2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n881), .A3(new_n312), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n858), .A2(new_n861), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n850), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n312), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n883), .B1(new_n888), .B2(G148gat), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n859), .A2(new_n862), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT59), .B(new_n881), .C1(new_n890), .C2(new_n312), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n882), .B1(new_n889), .B2(new_n891), .ZN(G1345gat));
  INV_X1    g691(.A(G155gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n893), .A3(new_n289), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n890), .A2(new_n289), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n893), .ZN(G1346gat));
  NAND2_X1  g695(.A1(new_n890), .A2(new_n693), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G162gat), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n265), .A2(G162gat), .A3(new_n553), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n866), .B2(new_n899), .ZN(G1347gat));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n651), .A2(new_n554), .ZN(new_n902));
  INV_X1    g701(.A(new_n842), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n860), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT121), .B(new_n904), .C1(new_n832), .C2(new_n833), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n340), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n904), .B1(new_n832), .B2(new_n833), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT119), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n376), .A3(new_n737), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(G1348gat));
  NAND3_X1  g716(.A1(new_n908), .A2(G176gat), .A3(new_n312), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  AOI21_X1  g720(.A(G176gat), .B1(new_n912), .B2(new_n312), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(G1349gat));
  AND3_X1   g722(.A1(new_n911), .A2(new_n384), .A3(new_n289), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n289), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(G183gat), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1350gat));
  AOI21_X1  g727(.A(new_n385), .B1(new_n908), .B2(new_n693), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT124), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n860), .A2(new_n905), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n911), .A2(new_n901), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n693), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G190gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n930), .A3(G190gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n935), .A2(KEYINPUT125), .A3(new_n930), .A4(G190gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n931), .A2(new_n938), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n912), .A2(new_n385), .A3(new_n693), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1351gat));
  NAND4_X1  g744(.A1(new_n672), .A2(new_n521), .A3(new_n599), .A4(new_n553), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n832), .B2(new_n833), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n737), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n672), .A2(new_n902), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n886), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n737), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  NAND3_X1  g752(.A1(new_n886), .A2(new_n312), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n947), .A2(new_n956), .A3(new_n312), .ZN(new_n957));
  OR3_X1    g756(.A1(new_n957), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT126), .B1(new_n957), .B2(KEYINPUT62), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n958), .A2(new_n959), .B1(KEYINPUT62), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n955), .A2(new_n960), .ZN(G1353gat));
  INV_X1    g760(.A(G211gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n962), .A3(new_n289), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n289), .B(new_n950), .C1(new_n884), .C2(new_n885), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n947), .B2(new_n693), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT127), .Z(new_n969));
  AND2_X1   g768(.A1(new_n693), .A2(G218gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n951), .B2(new_n970), .ZN(G1355gat));
endmodule


