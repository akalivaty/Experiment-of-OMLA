//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT66), .Z(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n466), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n464), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n467), .A2(new_n469), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n489), .B(new_n490), .C1(new_n465), .C2(new_n466), .ZN(new_n491));
  AND2_X1   g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n469), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n480), .B2(new_n490), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n465), .B2(new_n466), .ZN(new_n496));
  AND2_X1   g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n503), .A2(new_n505), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n511), .A2(new_n513), .A3(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n509), .A2(new_n516), .A3(new_n519), .A4(KEYINPUT68), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G62), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n510), .B1(new_n523), .B2(new_n501), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n514), .A2(new_n525), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n521), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(new_n528), .ZN(G166));
  AOI22_X1  g104(.A1(new_n515), .A2(G89), .B1(new_n518), .B2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G168));
  XOR2_X1   g111(.A(KEYINPUT71), .B(G90), .Z(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n514), .A2(new_n537), .B1(new_n517), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT6), .B(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT71), .B(G90), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n522), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n549), .A2(new_n542), .A3(G543), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n544), .A2(new_n550), .A3(KEYINPUT72), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n541), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n522), .A2(G64), .ZN(new_n553));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n510), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT73), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  AOI211_X1 g133(.A(new_n558), .B(new_n555), .C1(new_n541), .C2(new_n551), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  AOI22_X1  g136(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(new_n510), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT75), .B(G81), .Z(new_n564));
  XOR2_X1   g139(.A(KEYINPUT74), .B(G43), .Z(new_n565));
  OAI22_X1  g140(.A1(new_n514), .A2(new_n564), .B1(new_n565), .B2(new_n517), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n503), .A2(new_n505), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n503), .B2(new_n505), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n579), .B2(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n580), .B2(new_n510), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n522), .A2(new_n576), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n582), .A2(new_n583), .A3(G65), .ZN(new_n584));
  INV_X1    g159(.A(new_n575), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(G651), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n542), .A2(KEYINPUT76), .A3(G543), .ZN(new_n589));
  INV_X1    g164(.A(G53), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT9), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT9), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n592), .A4(G53), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n591), .A2(new_n593), .B1(G91), .B2(new_n515), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n581), .A2(new_n588), .A3(new_n594), .ZN(G299));
  INV_X1    g170(.A(G168), .ZN(G286));
  INV_X1    g171(.A(G166), .ZN(G303));
  NAND2_X1  g172(.A1(new_n515), .A2(G87), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n518), .A2(G49), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G288));
  AOI22_X1  g176(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n510), .ZN(new_n603));
  INV_X1    g178(.A(G86), .ZN(new_n604));
  INV_X1    g179(.A(G48), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n514), .A2(new_n604), .B1(new_n517), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n603), .A2(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n510), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n514), .A2(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND3_X1  g189(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n514), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n518), .A2(G54), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n579), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n510), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G171), .B2(new_n623), .ZN(G284));
  OAI21_X1  g200(.A(new_n624), .B1(G171), .B2(new_n623), .ZN(G321));
  NAND2_X1  g201(.A1(G299), .A2(new_n623), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n623), .B2(G168), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n623), .B2(G168), .ZN(G280));
  INV_X1    g204(.A(new_n622), .ZN(new_n630));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n481), .A2(G2104), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n481), .A2(G135), .ZN(new_n641));
  OR2_X1    g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(G123), .B2(new_n483), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n640), .A2(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(KEYINPUT81), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT80), .B(KEYINPUT14), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n663), .A3(new_n661), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n669), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n670), .ZN(new_n676));
  INV_X1    g251(.A(new_n669), .ZN(new_n677));
  OR3_X1    g252(.A1(new_n672), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n669), .A3(new_n670), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT84), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n684), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n694), .B1(KEYINPUT20), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n697), .B(new_n698), .C1(KEYINPUT20), .C2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT85), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n704), .A2(new_n705), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  NOR2_X1   g284(.A1(G16), .A2(G21), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G168), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1966), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G33), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G103), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n481), .A2(G139), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n717), .B(new_n718), .C1(new_n469), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n712), .B1(G2072), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT98), .B(KEYINPUT30), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G28), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(new_n713), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n645), .B2(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n722), .B2(G2072), .ZN(new_n728));
  NOR2_X1   g303(.A1(G164), .A2(new_n713), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G27), .B2(new_n713), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n728), .B1(G2078), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(G29), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n481), .A2(G141), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT96), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n483), .A2(G129), .B1(G105), .B2(new_n476), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(new_n713), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n734), .B(new_n744), .C1(new_n742), .C2(new_n713), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n733), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT97), .B(KEYINPUT31), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G11), .ZN(new_n753));
  NOR2_X1   g328(.A1(G5), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G171), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1961), .Z(new_n756));
  AND2_X1   g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  NOR2_X1   g332(.A1(KEYINPUT24), .A2(G34), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n757), .A2(new_n758), .A3(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n478), .B2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT95), .B(G2084), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n751), .A2(new_n753), .A3(new_n756), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G20), .ZN(new_n770));
  MUX2_X1   g345(.A(new_n767), .B(new_n768), .S(new_n770), .Z(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n630), .B2(new_n769), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(G1348), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n775), .B(new_n776), .Z(new_n777));
  AND2_X1   g352(.A1(new_n713), .A2(G26), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n481), .A2(G140), .B1(G128), .B2(new_n483), .ZN(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT92), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n464), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n782), .B1(new_n781), .B2(new_n780), .C1(G116), .C2(new_n469), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(G29), .ZN(new_n785));
  MUX2_X1   g360(.A(new_n778), .B(new_n785), .S(KEYINPUT28), .Z(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT93), .B(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n769), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n567), .B2(new_n769), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1341), .Z(new_n791));
  NAND4_X1  g366(.A1(new_n773), .A2(new_n777), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n771), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(G1956), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n765), .A2(new_n766), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n769), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(G288), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n769), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT33), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1976), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n769), .A2(G6), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n603), .A2(new_n606), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n769), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT89), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G22), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G166), .B2(G16), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1971), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n800), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n769), .A2(G24), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n613), .B2(new_n769), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n818));
  INV_X1    g393(.A(G95), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n469), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT87), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n483), .A2(G119), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n481), .A2(G131), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  INV_X1    g400(.A(G25), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT86), .B1(new_n826), .B2(G29), .ZN(new_n827));
  OR3_X1    g402(.A1(new_n826), .A2(KEYINPUT86), .A3(G29), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT35), .B(G1991), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n810), .A2(new_n812), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n813), .A2(new_n817), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n713), .A2(G35), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G162), .B2(new_n713), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT29), .B(G2090), .Z(new_n840));
  XOR2_X1   g415(.A(new_n839), .B(new_n840), .Z(new_n841));
  NOR4_X1   g416(.A1(new_n795), .A2(new_n836), .A3(new_n837), .A4(new_n841), .ZN(G311));
  INV_X1    g417(.A(G311), .ZN(G150));
  XNOR2_X1  g418(.A(KEYINPUT102), .B(G93), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n515), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n518), .A2(G55), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n503), .A2(new_n505), .A3(G67), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n847), .B1(new_n850), .B2(G651), .ZN(new_n851));
  AOI211_X1 g426(.A(KEYINPUT101), .B(new_n510), .C1(new_n848), .C2(new_n849), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n845), .B(new_n846), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n622), .A2(new_n631), .ZN(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT39), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n563), .A2(new_n566), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n853), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n855), .B1(new_n862), .B2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT103), .Z(G145));
  NAND2_X1  g439(.A1(new_n499), .A2(KEYINPUT104), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n493), .A2(new_n866), .A3(new_n494), .A4(new_n498), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n784), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n720), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n638), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n481), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n483), .A2(G130), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n869), .B(new_n720), .ZN(new_n878));
  INV_X1    g453(.A(new_n638), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n871), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n877), .B1(new_n871), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n742), .B(new_n824), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n645), .B(new_n487), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n886), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(G160), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G160), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT105), .B(G37), .Z(new_n893));
  OAI22_X1  g468(.A1(new_n881), .A2(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  AND3_X1   g471(.A1(new_n520), .A2(new_n528), .A3(G288), .ZN(new_n897));
  AOI21_X1  g472(.A(G288), .B1(new_n520), .B2(new_n528), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n802), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(G166), .A2(new_n797), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n520), .A2(new_n528), .A3(G288), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(G305), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n899), .A2(new_n902), .A3(new_n613), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n613), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n587), .B1(new_n586), .B2(G651), .ZN(new_n908));
  AOI211_X1 g483(.A(KEYINPUT79), .B(new_n510), .C1(new_n584), .C2(new_n585), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n594), .A3(new_n622), .ZN(new_n911));
  NAND2_X1  g486(.A1(G299), .A2(new_n630), .ZN(new_n912));
  AOI211_X1 g487(.A(new_n907), .B(KEYINPUT41), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT41), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT41), .B1(new_n911), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n861), .B(new_n633), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n911), .A2(new_n912), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n918), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n906), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n917), .A2(new_n918), .ZN(new_n924));
  INV_X1    g499(.A(new_n922), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT42), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n905), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(new_n906), .A3(new_n922), .ZN(new_n928));
  INV_X1    g503(.A(new_n905), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n924), .B2(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n623), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n853), .A2(new_n623), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n923), .A2(new_n926), .A3(new_n905), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(G295));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n933), .ZN(G331));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n853), .B(new_n567), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n544), .A2(new_n550), .A3(KEYINPUT72), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT72), .B1(new_n544), .B2(new_n550), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n556), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n558), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n552), .A2(KEYINPUT73), .A3(new_n556), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n949), .A2(G168), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G286), .B1(new_n557), .B2(new_n559), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(new_n950), .A3(G168), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n861), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(KEYINPUT109), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n954), .A2(new_n861), .A3(new_n958), .A4(new_n955), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n961), .A3(new_n956), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(new_n861), .A3(KEYINPUT110), .A4(new_n955), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n917), .A2(new_n960), .B1(new_n920), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n903), .B2(new_n904), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n899), .A2(new_n902), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G290), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n899), .A2(new_n902), .A3(new_n613), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(KEYINPUT111), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n943), .B(new_n944), .C1(new_n965), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(new_n920), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT41), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n920), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT41), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n907), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n915), .A2(KEYINPUT107), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n957), .A3(new_n979), .A4(new_n959), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n972), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT112), .B1(new_n981), .B2(G37), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n965), .A2(new_n905), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n973), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n972), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n960), .A2(new_n921), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n964), .A2(new_n916), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n983), .A2(new_n990), .A3(new_n893), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n985), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(G397));
  INV_X1    g575(.A(new_n742), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n784), .B(G2067), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n742), .A2(G1996), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n824), .A2(new_n830), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT124), .ZN(new_n1008));
  OAI22_X1  g583(.A1(new_n1006), .A2(new_n1008), .B1(G2067), .B2(new_n784), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n865), .B2(new_n867), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT45), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n470), .A2(new_n475), .A3(G40), .A4(new_n477), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT125), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(KEYINPUT46), .A3(new_n1002), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n1014), .B2(G1996), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1018), .B(new_n1020), .C1(new_n1014), .C2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  INV_X1    g598(.A(new_n1006), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n824), .A2(new_n830), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1007), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1015), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT126), .Z(new_n1028));
  NAND3_X1  g603(.A1(new_n1015), .A2(new_n816), .A3(new_n613), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1017), .B(new_n1023), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT55), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n499), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1012), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n1037), .B(G1384), .C1(new_n865), .C2(new_n867), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT113), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1010), .A2(KEYINPUT45), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1038), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n1035), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT50), .B1(new_n499), .B2(new_n1035), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1013), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(G8), .B(new_n1034), .C1(new_n1045), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1036), .A2(new_n1012), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n802), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(new_n1062), .A3(new_n1058), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1060), .A2(KEYINPUT116), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1055), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT117), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n797), .A2(G1976), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1054), .A2(G8), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(KEYINPUT114), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1072), .B(new_n1074), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n797), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1068), .A2(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1053), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1058), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1976), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(new_n797), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1081), .B2(new_n1055), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1036), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1012), .B1(new_n1084), .B2(new_n1046), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(G1961), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1038), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1087), .A2(new_n1088), .A3(G2078), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1041), .A2(new_n747), .A3(new_n1044), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(KEYINPUT123), .A3(new_n1092), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1086), .B(new_n1089), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(G8), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1033), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1077), .A3(new_n1052), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G286), .A2(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT121), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT51), .ZN(new_n1104));
  INV_X1    g679(.A(G1966), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1087), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2084), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1085), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(new_n1104), .C1(new_n1109), .C2(G286), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(G8), .A3(G286), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1104), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1087), .A2(new_n1105), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1113));
  INV_X1    g688(.A(G8), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(new_n1102), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1110), .A2(new_n1115), .A3(KEYINPUT62), .A4(new_n1111), .ZN(new_n1119));
  AOI21_X1  g694(.A(G301), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1082), .B1(new_n1101), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1042), .A2(new_n1038), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1049), .A2(new_n772), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT57), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(KEYINPUT57), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(G299), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OR3_X1    g704(.A1(G299), .A2(new_n1125), .A3(KEYINPUT57), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1123), .A2(new_n1124), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1123), .A2(new_n1124), .B1(new_n1130), .B2(new_n1129), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1085), .A2(new_n776), .B1(new_n1054), .B2(G2067), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT119), .A3(new_n630), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT119), .B1(new_n1134), .B2(new_n630), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1131), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(new_n630), .ZN(new_n1139));
  OAI221_X1 g714(.A(new_n622), .B1(new_n1054), .B2(G2067), .C1(new_n1085), .C2(new_n776), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT120), .B(G1996), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1042), .A2(new_n1038), .A3(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  AND2_X1   g719(.A1(new_n1054), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n567), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1141), .A2(KEYINPUT60), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1131), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1132), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1133), .A2(KEYINPUT61), .A3(new_n1131), .ZN(new_n1152));
  OR3_X1    g727(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n622), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1138), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G301), .B(KEYINPUT54), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1086), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1096), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1157), .B1(new_n1161), .B2(new_n1089), .ZN(new_n1162));
  AND4_X1   g737(.A1(new_n1116), .A2(new_n1099), .A3(new_n1077), .A4(new_n1052), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1011), .A2(new_n1040), .A3(new_n1012), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1088), .A2(G2078), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1157), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1158), .B(new_n1166), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1113), .A2(new_n1114), .A3(G286), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1099), .A2(new_n1077), .A3(new_n1052), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1121), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1026), .B1(G1986), .B2(G290), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(G1986), .B2(G290), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1175), .A2(new_n1015), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1031), .B1(new_n1173), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g752(.A1(new_n687), .A2(new_n667), .ZN(new_n1179));
  INV_X1    g753(.A(new_n461), .ZN(new_n1180));
  OAI21_X1  g754(.A(new_n1180), .B1(new_n707), .B2(new_n708), .ZN(new_n1181));
  OAI21_X1  g755(.A(KEYINPUT127), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(new_n708), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n461), .B1(new_n1183), .B2(new_n706), .ZN(new_n1184));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1185));
  NAND4_X1  g759(.A1(new_n1184), .A2(new_n1185), .A3(new_n667), .A4(new_n687), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n997), .A2(new_n1187), .A3(new_n895), .ZN(G225));
  INV_X1    g762(.A(G225), .ZN(G308));
endmodule


