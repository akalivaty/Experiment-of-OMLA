//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G50), .A2(G226), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n210), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT65), .Z(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n215), .B(new_n229), .C1(new_n231), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n230), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n209), .B2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n202), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n260), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(G20), .B2(new_n203), .ZN(new_n268));
  INV_X1    g0068(.A(new_n254), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n256), .B(new_n259), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  OAI211_X1 g0072(.A(G1), .B(G13), .C1(new_n261), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G1698), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G222), .B2(G1698), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G77), .B2(new_n277), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n272), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n209), .A4(G274), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n230), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n272), .B2(new_n284), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G226), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n279), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G200), .B2(new_n293), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n271), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT69), .B1(new_n293), .B2(G200), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n297), .B(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n293), .A2(G179), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n270), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n274), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n277), .B(new_n308), .C1(G226), .C2(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n289), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n273), .A2(G232), .A3(new_n281), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n287), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n303), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n273), .B1(new_n309), .B2(new_n310), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n317), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n265), .A2(G159), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT75), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n225), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n325), .B2(new_n201), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n328), .B(G20), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT74), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n329), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n329), .B2(new_n331), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n210), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n336), .B2(new_n328), .ZN(new_n337));
  OAI211_X1 g0137(.A(KEYINPUT16), .B(new_n327), .C1(new_n337), .C2(new_n225), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n323), .A2(new_n326), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n328), .B1(new_n277), .B2(G20), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n329), .A2(new_n331), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n225), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(new_n254), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n260), .A2(new_n257), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n255), .B2(new_n260), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT76), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n320), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT18), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n312), .A2(G190), .A3(new_n315), .ZN(new_n352));
  OAI21_X1  g0152(.A(G200), .B1(new_n317), .B2(new_n314), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n346), .A2(new_n352), .A3(new_n349), .A4(new_n353), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT17), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(KEYINPUT77), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n255), .A2(G77), .ZN(new_n361));
  XOR2_X1   g0161(.A(new_n361), .B(KEYINPUT68), .Z(new_n362));
  INV_X1    g0162(.A(new_n260), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n364));
  XOR2_X1   g0164(.A(KEYINPUT15), .B(G87), .Z(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n262), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n367), .A2(new_n269), .B1(G77), .B2(new_n257), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n277), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n342), .A2(new_n237), .A3(G1698), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n289), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n291), .A2(G244), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n287), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n303), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n377), .A2(G179), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(G200), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n369), .B(new_n381), .C1(new_n294), .C2(new_n377), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n306), .A2(new_n360), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n283), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT70), .B1(new_n283), .B2(new_n286), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n291), .A2(G238), .ZN(new_n389));
  INV_X1    g0189(.A(G97), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n261), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G226), .A2(G1698), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n237), .B2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n393), .B2(new_n277), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n389), .B1(new_n273), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT13), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n237), .A2(G1698), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G226), .B2(G1698), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n398), .A2(new_n342), .B1(new_n261), .B2(new_n390), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n289), .B1(G238), .B2(new_n291), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n387), .C2(new_n386), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(KEYINPUT13), .C1(new_n388), .C2(new_n395), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G179), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n396), .A2(new_n402), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n303), .B1(new_n396), .B2(new_n402), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT14), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n255), .A2(G68), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n258), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT12), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n257), .B2(G68), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT72), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n262), .A2(G77), .B1(G20), .B2(new_n225), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n265), .A2(G50), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n269), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g0224(.A(new_n424), .B(KEYINPUT11), .Z(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n408), .A2(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(new_n406), .B2(G190), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n414), .A2(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n384), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n209), .A2(G33), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n269), .A2(new_n434), .A3(new_n257), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n390), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n257), .A2(G97), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT7), .B1(new_n342), .B2(new_n210), .ZN(new_n438));
  OAI21_X1  g0238(.A(G107), .B1(new_n438), .B2(new_n332), .ZN(new_n439));
  INV_X1    g0239(.A(G77), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT78), .B1(new_n266), .B2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n266), .A2(KEYINPUT78), .A3(new_n440), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT6), .ZN(new_n443));
  AND2_X1   g0243(.A1(G97), .A2(G107), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n206), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n372), .A2(KEYINPUT6), .A3(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n442), .B1(new_n447), .B2(G20), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n439), .A2(new_n441), .A3(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n436), .B(new_n437), .C1(new_n449), .C2(new_n254), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G41), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n209), .B(G45), .C1(new_n272), .C2(KEYINPUT5), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n273), .B(new_n453), .C1(new_n454), .C2(KEYINPUT80), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n282), .B1(new_n454), .B2(KEYINPUT80), .ZN(new_n457));
  INV_X1    g0257(.A(new_n454), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n289), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(G257), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n329), .A2(new_n331), .A3(G244), .A4(new_n307), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT4), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n329), .A2(new_n331), .A3(G250), .A4(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n460), .B1(new_n469), .B2(new_n273), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G200), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n460), .B(G190), .C1(new_n469), .C2(new_n273), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n450), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n449), .A2(new_n254), .ZN(new_n474));
  INV_X1    g0274(.A(new_n436), .ZN(new_n475));
  INV_X1    g0275(.A(new_n437), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n303), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n460), .B(new_n318), .C1(new_n469), .C2(new_n273), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n365), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n258), .ZN(new_n483));
  INV_X1    g0283(.A(new_n435), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n365), .ZN(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(new_n391), .B2(KEYINPUT19), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT82), .B(G87), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT83), .B1(new_n487), .B2(new_n207), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n217), .A2(KEYINPUT82), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(new_n206), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n486), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n342), .A2(G20), .A3(new_n225), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT19), .B1(new_n262), .B2(G97), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n483), .B(new_n485), .C1(new_n498), .C2(new_n269), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n209), .A2(G45), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(G250), .C1(new_n288), .C2(new_n230), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n226), .A2(new_n307), .ZN(new_n503));
  INV_X1    g0303(.A(G244), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G1698), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n329), .A2(new_n503), .A3(new_n331), .A4(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n509), .B2(new_n289), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n500), .A2(new_n282), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G169), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n273), .B1(new_n506), .B2(new_n508), .ZN(new_n514));
  NOR4_X1   g0314(.A1(new_n514), .A2(G179), .A3(new_n502), .A4(new_n511), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT81), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n499), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n509), .A2(new_n289), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n294), .A3(new_n512), .A4(new_n501), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n514), .A2(new_n511), .A3(new_n502), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(new_n486), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n487), .A2(KEYINPUT83), .A3(new_n207), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n493), .B1(new_n492), .B2(new_n206), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n496), .ZN(new_n527));
  INV_X1    g0327(.A(new_n497), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n254), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n484), .A2(G87), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n522), .A2(new_n530), .A3(new_n531), .A4(new_n483), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n518), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n481), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n330), .A2(G33), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n536));
  OAI21_X1  g0336(.A(G303), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n329), .A2(new_n331), .A3(G257), .A4(new_n307), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n329), .A2(new_n331), .A3(G264), .A4(G1698), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT84), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n289), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(G270), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n303), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n484), .A2(G116), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n258), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n253), .A2(new_n230), .B1(G20), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n467), .B(new_n210), .C1(G33), .C2(new_n390), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT20), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n550), .A2(KEYINPUT20), .A3(new_n551), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n547), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n546), .A2(KEYINPUT21), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT21), .B1(new_n546), .B2(new_n554), .ZN(new_n556));
  INV_X1    g0356(.A(new_n554), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n544), .A2(new_n545), .A3(G179), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n544), .A2(new_n545), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(new_n557), .C1(new_n294), .C2(new_n561), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n534), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n435), .A2(new_n372), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n210), .B2(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(new_n210), .B2(new_n507), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n567), .B(KEYINPUT23), .C1(new_n210), .C2(G107), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n329), .A2(new_n331), .A3(new_n210), .A4(G87), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT85), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT24), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n568), .A2(new_n569), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n507), .A2(new_n210), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(new_n571), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n573), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(new_n210), .A3(G87), .A4(new_n277), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n581), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n254), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT87), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n590), .A3(new_n254), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n566), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n257), .A2(G107), .ZN(new_n593));
  XNOR2_X1  g0393(.A(new_n593), .B(KEYINPUT25), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n273), .B(G264), .C1(new_n454), .C2(new_n452), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n329), .A2(new_n331), .A3(G250), .A4(new_n307), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT88), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT88), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n277), .A2(new_n599), .A3(G250), .A4(new_n307), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G294), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n277), .A2(G257), .A3(G1698), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n596), .B1(new_n603), .B2(new_n289), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n456), .A2(new_n457), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G200), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(G190), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n592), .A2(new_n594), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  INV_X1    g0413(.A(new_n566), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n590), .B1(new_n587), .B2(new_n254), .ZN(new_n615));
  AOI211_X1 g0415(.A(KEYINPUT87), .B(new_n269), .C1(new_n578), .C2(new_n586), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n594), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(G169), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n318), .B2(new_n606), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n612), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n613), .B1(new_n612), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n565), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n433), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n305), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n428), .A2(new_n427), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n411), .B(KEYINPUT14), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(new_n407), .B1(new_n421), .B2(new_n425), .ZN(new_n628));
  INV_X1    g0428(.A(new_n380), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n359), .B(new_n626), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n351), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n625), .B1(new_n631), .B2(new_n301), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n620), .A2(new_n560), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n513), .A2(new_n515), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n499), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n473), .A2(new_n480), .A3(new_n532), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n617), .A2(new_n609), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n611), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n620), .A2(new_n560), .A3(KEYINPUT90), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  INV_X1    g0443(.A(new_n637), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n532), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n480), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n518), .A2(new_n532), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n649), .B2(new_n480), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(new_n647), .A3(new_n532), .A4(new_n637), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n650), .A2(new_n653), .A3(new_n643), .A4(new_n637), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n642), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n632), .B1(new_n433), .B2(new_n657), .ZN(G369));
  INV_X1    g0458(.A(G13), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G20), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n209), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n617), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n621), .B2(new_n622), .ZN(new_n668));
  INV_X1    g0468(.A(new_n666), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n620), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n560), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n557), .A2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n564), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n620), .A2(new_n666), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n560), .A2(new_n666), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n672), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n680), .A2(new_n684), .ZN(G399));
  NOR2_X1   g0485(.A1(new_n524), .A2(new_n525), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n548), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n213), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n232), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT95), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n696), .C1(new_n657), .C2(new_n666), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n647), .B1(new_n533), .B2(new_n652), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n437), .B1(new_n449), .B2(new_n254), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n699), .A2(new_n475), .B1(new_n470), .B2(new_n303), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n637), .A3(new_n479), .A4(new_n532), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n637), .B1(new_n701), .B2(KEYINPUT26), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT91), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n654), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n666), .B1(new_n704), .B2(new_n642), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT95), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n533), .A2(new_n647), .A3(new_n652), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n644), .B1(new_n701), .B2(KEYINPUT26), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n640), .B1(KEYINPUT96), .B2(new_n633), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n707), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .A3(new_n669), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n697), .A2(new_n706), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G330), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n565), .B(new_n669), .C1(new_n621), .C2(new_n622), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n604), .A2(new_n521), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n558), .A2(new_n470), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT30), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n558), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n459), .A2(G257), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n605), .A2(new_n721), .ZN(new_n722));
  OR3_X1    g0522(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n289), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n720), .A2(new_n604), .A3(new_n724), .A4(new_n521), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(KEYINPUT94), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n607), .A2(new_n724), .ZN(new_n728));
  INV_X1    g0528(.A(new_n521), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n728), .A2(new_n318), .A3(new_n561), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n719), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n666), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n731), .B2(new_n666), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n714), .B1(new_n715), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n713), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n694), .B1(new_n738), .B2(G1), .ZN(G364));
  AOI21_X1  g0539(.A(new_n230), .B1(G20), .B2(new_n303), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n210), .A2(new_n294), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n318), .A2(new_n608), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n210), .A2(G190), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n318), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n743), .A2(new_n202), .B1(new_n746), .B2(new_n440), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n741), .A2(new_n745), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(G58), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT98), .Z(new_n751));
  NOR2_X1   g0551(.A1(new_n608), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT99), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n372), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n741), .A2(new_n752), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n210), .B1(new_n758), .B2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(new_n487), .B1(new_n760), .B2(G97), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n742), .A2(new_n744), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n761), .B(new_n277), .C1(new_n225), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n758), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT32), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n751), .A2(new_n755), .A3(new_n763), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n277), .B1(new_n760), .B2(G294), .ZN(new_n771));
  INV_X1    g0571(.A(G303), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n771), .B1(new_n772), .B2(new_n756), .C1(new_n773), .C2(new_n746), .ZN(new_n774));
  INV_X1    g0574(.A(G326), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n743), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n762), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n765), .A2(G329), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n749), .A2(G322), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n770), .A2(new_n774), .A3(new_n776), .A4(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n740), .B1(new_n768), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n213), .A2(G355), .A3(new_n277), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n248), .A2(new_n284), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT74), .B1(new_n535), .B2(new_n536), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n329), .A2(new_n331), .A3(new_n333), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n689), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n233), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n787), .B1(G116), .B2(new_n213), .C1(new_n788), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n740), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n660), .A2(G45), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n691), .A2(G1), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n786), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  INV_X1    g0605(.A(new_n798), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n677), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n677), .A2(G330), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n678), .A2(new_n802), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n370), .A2(new_n666), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n380), .A2(new_n382), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n380), .A2(new_n811), .A3(new_n382), .A4(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n656), .A2(new_n669), .A3(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n814), .A2(new_n815), .B1(new_n629), .B2(new_n666), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n818), .B1(new_n705), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(new_n736), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n736), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n802), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n754), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n277), .B1(new_n825), .B2(G87), .ZN(new_n826));
  INV_X1    g0626(.A(new_n743), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G303), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n757), .A2(G107), .B1(new_n760), .B2(G97), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n762), .A2(new_n769), .B1(new_n746), .B2(new_n548), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n748), .A2(new_n831), .B1(new_n764), .B2(new_n773), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n826), .A2(new_n828), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G143), .A2(new_n749), .B1(new_n777), .B2(G150), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(G159), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n743), .C1(new_n837), .C2(new_n746), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n791), .B(new_n840), .C1(G50), .C2(new_n757), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n839), .A2(KEYINPUT34), .B1(G68), .B2(new_n825), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(new_n324), .C2(new_n759), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n764), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n834), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n740), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n740), .A2(new_n796), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n440), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n819), .A2(new_n796), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n803), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n824), .A2(new_n851), .ZN(G384));
  NAND2_X1  g0652(.A1(new_n432), .A2(new_n735), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n426), .A2(new_n666), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n429), .A2(new_n854), .B1(new_n628), .B2(new_n666), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n819), .B(new_n855), .C1(new_n715), .C2(new_n734), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n338), .A2(new_n254), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT7), .B1(new_n791), .B2(new_n210), .ZN(new_n858));
  OAI21_X1  g0658(.A(G68), .B1(new_n858), .B2(new_n332), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n859), .B2(new_n327), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n349), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n664), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT103), .B(new_n349), .C1(new_n857), .C2(new_n860), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n320), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n863), .A2(new_n867), .A3(new_n865), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n868), .A3(new_n354), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n346), .A2(new_n349), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n867), .B2(new_n864), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n354), .ZN(new_n873));
  XNOR2_X1  g0673(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n866), .B1(new_n351), .B2(new_n359), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n875), .B1(new_n869), .B2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(new_n878), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n856), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XOR2_X1   g0686(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n887));
  NAND2_X1  g0687(.A1(new_n871), .A2(new_n864), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n351), .B2(new_n359), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n346), .A2(new_n349), .B1(new_n320), .B2(new_n664), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n874), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n873), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n872), .A2(new_n891), .A3(new_n354), .A4(new_n874), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n887), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT107), .B(new_n887), .C1(new_n889), .C2(new_n895), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n880), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n885), .B1(new_n900), .B2(new_n856), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n886), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n853), .B1(new_n902), .B2(new_n714), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n856), .A2(new_n884), .A3(new_n885), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n900), .A2(new_n856), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n905), .B2(new_n885), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n715), .A2(new_n734), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n432), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n697), .A2(new_n706), .A3(new_n432), .A4(new_n712), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n632), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n884), .A2(KEYINPUT39), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n880), .A2(new_n898), .A3(new_n914), .A4(new_n899), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(KEYINPUT108), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n414), .A2(new_n426), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n666), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n898), .A2(new_n899), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT108), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n914), .A4(new_n880), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n916), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n666), .B(new_n816), .C1(new_n704), .C2(new_n642), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n380), .A2(new_n666), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n818), .A2(KEYINPUT102), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n855), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n884), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n351), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n664), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n922), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n912), .B(new_n934), .Z(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n209), .B2(new_n660), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n548), .B1(new_n447), .B2(KEYINPUT35), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(new_n231), .C1(KEYINPUT35), .C2(new_n447), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  OAI21_X1  g0739(.A(G77), .B1(new_n324), .B2(new_n225), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n940), .A2(new_n232), .B1(G50), .B2(new_n225), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n659), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n936), .A2(new_n939), .A3(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n481), .B1(new_n450), .B2(new_n669), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n652), .A2(new_n666), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n672), .A2(new_n682), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT42), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n480), .B1(new_n944), .B2(new_n620), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n669), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n530), .A2(new_n531), .A3(new_n483), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n666), .ZN(new_n955));
  MUX2_X1   g0755(.A(new_n637), .B(new_n645), .S(new_n955), .Z(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n953), .A2(KEYINPUT43), .A3(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n680), .A2(new_n946), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n958), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n959), .B1(new_n958), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n690), .B(KEYINPUT41), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n672), .A2(new_n682), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n672), .A2(new_n682), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT110), .B1(new_n677), .B2(G330), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n737), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT44), .B1(new_n683), .B2(new_n946), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n683), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n683), .A2(new_n946), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT45), .B1(new_n683), .B2(new_n946), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n979), .B(new_n980), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT109), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n986), .A3(new_n680), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n980), .A2(new_n979), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n981), .B(new_n982), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT109), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n978), .B(new_n987), .C1(new_n990), .C2(new_n680), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n968), .B1(new_n991), .B2(new_n738), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n801), .A2(G1), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n966), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G143), .A2(new_n827), .B1(new_n757), .B2(G58), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n440), .B2(new_n753), .C1(new_n836), .C2(new_n764), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n277), .B1(new_n759), .B2(new_n225), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n264), .A2(new_n748), .B1(new_n762), .B2(new_n837), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n202), .B2(new_n746), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n743), .A2(new_n773), .B1(new_n753), .B2(new_n390), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n756), .A2(new_n548), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(KEYINPUT46), .B1(new_n769), .B2(new_n746), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(KEYINPUT46), .C2(new_n1002), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT111), .B(G317), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n764), .A2(new_n1005), .B1(new_n759), .B2(new_n372), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1006), .B(new_n792), .C1(G294), .C2(new_n777), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1004), .B(new_n1007), .C1(new_n772), .C2(new_n748), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1000), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n740), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n956), .A2(new_n798), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n793), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n799), .B1(new_n213), .B2(new_n482), .C1(new_n1013), .C2(new_n243), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n803), .A4(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT112), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n994), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT113), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n994), .A2(KEYINPUT113), .A3(new_n1016), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(G387));
  NAND2_X1  g0821(.A1(new_n977), .A2(new_n737), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n738), .A2(new_n976), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n690), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n792), .B1(new_n754), .B2(new_n390), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n746), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(G68), .B2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n482), .A2(new_n759), .B1(new_n260), .B2(new_n762), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n743), .A2(new_n837), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n756), .A2(new_n440), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n764), .A2(new_n264), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1027), .B(new_n1032), .C1(new_n202), .C2(new_n748), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT115), .Z(new_n1034));
  AOI22_X1  g0834(.A1(G311), .A2(new_n777), .B1(new_n1026), .B2(G303), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n748), .B2(new_n1005), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT116), .B(G322), .Z(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n827), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT48), .Z(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n769), .B2(new_n759), .C1(new_n831), .C2(new_n756), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT49), .Z(new_n1041));
  OAI221_X1 g0841(.A(new_n791), .B1(new_n548), .B2(new_n753), .C1(new_n775), .C2(new_n764), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n740), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n673), .A2(new_n798), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n363), .A2(new_n1046), .A3(new_n202), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n688), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n225), .A2(new_n440), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n363), .B2(new_n202), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1048), .A2(G45), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n240), .A2(G45), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT114), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n793), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n687), .A2(new_n213), .A3(new_n277), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n213), .A2(G107), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n799), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1044), .A2(new_n803), .A3(new_n1045), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n993), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1024), .B(new_n1059), .C1(new_n1060), .C2(new_n977), .ZN(G393));
  AND2_X1   g0861(.A1(new_n985), .A2(new_n680), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n985), .A2(new_n680), .ZN(new_n1063));
  OR3_X1    g0863(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT117), .ZN(new_n1064));
  OAI21_X1  g0864(.A(KEYINPUT117), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n993), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1023), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n991), .A3(new_n690), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n944), .A2(new_n798), .A3(new_n945), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n799), .B1(new_n390), .B2(new_n213), .C1(new_n1013), .C2(new_n251), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n759), .A2(new_n440), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n792), .B1(new_n202), .B2(new_n762), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G143), .C2(new_n765), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1026), .A2(new_n363), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G150), .A2(new_n827), .B1(new_n749), .B2(G159), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n825), .A2(G87), .B1(KEYINPUT51), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(KEYINPUT51), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G68), .B2(new_n757), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G317), .A2(new_n827), .B1(new_n749), .B2(G311), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT52), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n342), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G283), .B2(new_n757), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1026), .A2(G294), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n755), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G303), .A2(new_n777), .B1(new_n765), .B2(new_n1037), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n759), .A2(new_n548), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1079), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n740), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1069), .A2(new_n803), .A3(new_n1070), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1066), .A2(new_n1068), .A3(new_n1092), .ZN(G390));
  NAND3_X1  g0893(.A1(new_n735), .A2(new_n820), .A3(new_n930), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n923), .B(new_n925), .C1(new_n705), .C2(new_n817), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT102), .B1(new_n818), .B2(new_n927), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n930), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n918), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1098), .A2(new_n1099), .B1(new_n916), .B2(new_n921), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n711), .A2(new_n669), .A3(new_n817), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n927), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1099), .B(new_n900), .C1(new_n1103), .C2(new_n855), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1095), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n918), .B1(new_n929), .B2(new_n930), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n915), .A2(KEYINPUT108), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n920), .B1(new_n884), .B2(KEYINPUT39), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n915), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1104), .B(new_n1094), .C1(new_n1107), .C2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1106), .A2(new_n1111), .A3(new_n993), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1110), .A2(new_n797), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n848), .A2(new_n260), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n762), .A2(new_n836), .B1(new_n764), .B2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  AOI211_X1 g0917(.A(new_n342), .B(new_n1116), .C1(new_n1026), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n760), .A2(G159), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT53), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n757), .A2(new_n1120), .A3(G150), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n757), .B2(G150), .ZN(new_n1122));
  INV_X1    g0922(.A(G128), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n743), .A2(new_n1123), .B1(new_n748), .B2(new_n844), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n753), .A2(new_n202), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .A4(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G107), .A2(new_n777), .B1(new_n1026), .B2(G97), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n825), .A2(G68), .B1(new_n1129), .B2(KEYINPUT118), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n277), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n748), .A2(new_n548), .B1(new_n764), .B2(new_n831), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1071), .B(new_n1133), .C1(G283), .C2(new_n827), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n756), .A2(new_n217), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1127), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n740), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1113), .A2(new_n803), .A3(new_n1114), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1112), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n910), .A2(new_n632), .A3(new_n853), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n930), .B1(new_n735), .B2(new_n820), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1095), .A2(new_n1142), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1103), .A2(new_n1144), .A3(new_n1094), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1141), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1106), .A2(new_n1111), .A3(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1147), .A2(new_n690), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1141), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1140), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(G378));
  XNOR2_X1  g0955(.A(new_n306), .B(KEYINPUT119), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n270), .A2(new_n864), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1156), .B(new_n1159), .Z(new_n1160));
  AOI21_X1  g0960(.A(new_n802), .B1(new_n1160), .B2(new_n796), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n482), .A2(new_n746), .B1(new_n390), .B2(new_n762), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1162), .A2(new_n792), .A3(G41), .A4(new_n1030), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n753), .A2(new_n324), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n748), .A2(new_n372), .B1(new_n764), .B2(new_n769), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G68), .C2(new_n760), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1163), .B(new_n1166), .C1(new_n548), .C2(new_n743), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT58), .Z(new_n1168));
  AOI21_X1  g0968(.A(G50), .B1(new_n791), .B2(new_n272), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(G33), .B2(G41), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G128), .A2(new_n749), .B1(new_n777), .B2(G132), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n827), .A2(G125), .B1(new_n760), .B2(G150), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n757), .A2(new_n1117), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1026), .A2(G137), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT59), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n837), .B2(new_n753), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1170), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n740), .B1(new_n1168), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n848), .A2(new_n202), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1161), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT120), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1160), .B1(new_n906), .B2(G330), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G330), .B(new_n1160), .C1(new_n886), .C2(new_n901), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n934), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1160), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n902), .B2(new_n714), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n855), .B1(new_n926), .B2(new_n928), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1190), .A2(new_n884), .B1(new_n932), .B2(new_n664), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n1191), .A3(new_n922), .A4(new_n1185), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1193), .B2(new_n1060), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1187), .A2(new_n1192), .A3(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n690), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1195), .B1(new_n1199), .B2(new_n1201), .ZN(G375));
  AOI22_X1  g1002(.A1(new_n825), .A2(G77), .B1(G294), .B2(new_n827), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n762), .A2(new_n548), .B1(new_n746), .B2(new_n372), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT121), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n277), .B1(new_n760), .B2(new_n365), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G283), .A2(new_n749), .B1(new_n765), .B2(G303), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G97), .B2(new_n757), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n756), .A2(new_n837), .B1(new_n764), .B2(new_n1123), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT122), .Z(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n792), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n748), .A2(new_n836), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1164), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n202), .B2(new_n759), .C1(new_n844), .C2(new_n743), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1117), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1216), .A2(new_n762), .B1(new_n746), .B2(new_n264), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n740), .B1(new_n1209), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n803), .B(new_n1219), .C1(new_n930), .C2(new_n797), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n225), .B2(new_n848), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1151), .B2(new_n993), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1141), .A2(new_n1145), .A3(new_n1143), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n967), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1224), .B2(new_n1146), .ZN(G381));
  INV_X1    g1025(.A(G390), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1019), .A2(new_n1020), .A3(new_n1226), .ZN(new_n1227));
  OR3_X1    g1027(.A1(new_n1227), .A2(G396), .A3(G393), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n691), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1194), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1154), .ZN(new_n1234));
  OR2_X1    g1034(.A1(G381), .A2(G384), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1228), .A2(new_n1234), .A3(new_n1235), .ZN(G407));
  OAI21_X1  g1036(.A(G343), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1154), .A3(new_n1233), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(G213), .ZN(G409));
  NAND3_X1  g1039(.A1(new_n1197), .A2(new_n1200), .A3(new_n967), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1154), .A2(new_n1195), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n665), .A2(G213), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n1233), .C2(new_n1154), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1223), .A2(KEYINPUT123), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n690), .B(new_n1152), .C1(new_n1244), .C2(KEYINPUT60), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(KEYINPUT60), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1222), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G384), .B(new_n1222), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n665), .A2(G213), .A3(G2897), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1243), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1255), .A2(new_n1256), .B1(new_n1243), .B2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(G393), .B(G396), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1017), .A2(G390), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1227), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1017), .B1(new_n1226), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1259), .B1(new_n1226), .B2(new_n1262), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(G390), .A2(new_n994), .A3(KEYINPUT124), .A4(new_n1016), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G375), .A2(G378), .B1(G213), .B2(new_n665), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1257), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(KEYINPUT63), .A3(new_n1241), .A4(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1258), .A2(new_n1268), .A3(new_n1269), .A4(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1270), .A2(new_n1274), .A3(new_n1241), .A4(new_n1271), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT62), .B1(new_n1243), .B2(new_n1257), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1243), .A2(new_n1254), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(new_n1269), .ZN(new_n1280));
  AOI211_X1 g1080(.A(KEYINPUT125), .B(KEYINPUT61), .C1(new_n1243), .C2(new_n1254), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1273), .B1(new_n1282), .B2(new_n1268), .ZN(G405));
  NAND2_X1  g1083(.A1(G375), .A2(G378), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1234), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1271), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1267), .A2(KEYINPUT126), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1261), .A2(new_n1288), .A3(new_n1266), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(G402));
endmodule


