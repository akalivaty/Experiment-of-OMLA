

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760;

  XOR2_X2 U361 ( .A(KEYINPUT69), .B(KEYINPUT0), .Z(n504) );
  INV_X1 U362 ( .A(G953), .ZN(n755) );
  AND2_X1 U363 ( .A1(n347), .A2(n345), .ZN(n340) );
  AND2_X2 U364 ( .A1(n392), .A2(n382), .ZN(n367) );
  XNOR2_X2 U365 ( .A(n376), .B(n535), .ZN(n644) );
  NOR2_X2 U366 ( .A1(n720), .A2(n716), .ZN(n569) );
  NAND2_X2 U367 ( .A1(n428), .A2(KEYINPUT2), .ZN(n427) );
  XOR2_X2 U368 ( .A(G137), .B(G131), .Z(n445) );
  NOR2_X2 U369 ( .A1(n556), .A2(n545), .ZN(n481) );
  NOR2_X1 U370 ( .A1(n346), .A2(n341), .ZN(n345) );
  NAND2_X1 U371 ( .A1(n340), .A2(n342), .ZN(n349) );
  AND2_X1 U372 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U373 ( .A1(n573), .A2(n574), .ZN(n418) );
  AND2_X1 U374 ( .A1(n429), .A2(KEYINPUT65), .ZN(n382) );
  NOR2_X1 U375 ( .A1(n550), .A2(n642), .ZN(n551) );
  NOR2_X1 U376 ( .A1(n622), .A2(G478), .ZN(n346) );
  AND2_X1 U377 ( .A1(n622), .A2(G478), .ZN(n348) );
  XNOR2_X1 U378 ( .A(n532), .B(n531), .ZN(n564) );
  INV_X1 U379 ( .A(n660), .ZN(n341) );
  XNOR2_X1 U380 ( .A(n486), .B(n461), .ZN(n744) );
  NAND2_X1 U381 ( .A1(n344), .A2(n343), .ZN(n342) );
  INV_X1 U382 ( .A(n622), .ZN(n343) );
  INV_X1 U383 ( .A(n362), .ZN(n344) );
  NAND2_X1 U384 ( .A1(n362), .A2(n348), .ZN(n347) );
  XNOR2_X1 U385 ( .A(n349), .B(n624), .ZN(G63) );
  XNOR2_X2 U386 ( .A(n351), .B(n350), .ZN(n436) );
  XNOR2_X2 U387 ( .A(G116), .B(KEYINPUT89), .ZN(n350) );
  XNOR2_X2 U388 ( .A(G119), .B(KEYINPUT3), .ZN(n351) );
  XNOR2_X2 U389 ( .A(n477), .B(n446), .ZN(n746) );
  NAND2_X1 U390 ( .A1(n368), .A2(n380), .ZN(n352) );
  BUF_X1 U391 ( .A(n743), .Z(n353) );
  NAND2_X1 U392 ( .A1(n368), .A2(n380), .ZN(n595) );
  XNOR2_X2 U393 ( .A(n483), .B(n482), .ZN(n736) );
  XNOR2_X2 U394 ( .A(n436), .B(n435), .ZN(n483) );
  NAND2_X1 U395 ( .A1(n410), .A2(KEYINPUT74), .ZN(n405) );
  INV_X1 U396 ( .A(n437), .ZN(n422) );
  OR2_X1 U397 ( .A1(n494), .A2(n490), .ZN(n440) );
  XNOR2_X1 U398 ( .A(n724), .B(KEYINPUT85), .ZN(n379) );
  INV_X1 U399 ( .A(KEYINPUT65), .ZN(n390) );
  AND2_X1 U400 ( .A1(n620), .A2(n390), .ZN(n389) );
  NOR2_X1 U401 ( .A1(n586), .A2(n587), .ZN(n601) );
  XNOR2_X1 U402 ( .A(n530), .B(G475), .ZN(n531) );
  NOR2_X1 U403 ( .A1(G902), .A2(n657), .ZN(n532) );
  INV_X1 U404 ( .A(KEYINPUT86), .ZN(n552) );
  INV_X1 U405 ( .A(n643), .ZN(n408) );
  XNOR2_X1 U406 ( .A(n606), .B(KEYINPUT47), .ZN(n410) );
  INV_X1 U407 ( .A(G237), .ZN(n491) );
  NOR2_X1 U408 ( .A1(G953), .A2(G237), .ZN(n521) );
  INV_X1 U409 ( .A(KEYINPUT4), .ZN(n370) );
  XNOR2_X1 U410 ( .A(G113), .B(KEYINPUT72), .ZN(n435) );
  XNOR2_X1 U411 ( .A(n414), .B(n413), .ZN(n507) );
  INV_X1 U412 ( .A(KEYINPUT8), .ZN(n413) );
  NAND2_X1 U413 ( .A1(n755), .A2(G234), .ZN(n414) );
  XNOR2_X1 U414 ( .A(G107), .B(G122), .ZN(n510) );
  XOR2_X1 U415 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n511) );
  XOR2_X1 U416 ( .A(G131), .B(G113), .Z(n519) );
  XNOR2_X1 U417 ( .A(G143), .B(G104), .ZN(n518) );
  XNOR2_X1 U418 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n485) );
  NAND2_X1 U419 ( .A1(G237), .A2(G234), .ZN(n498) );
  INV_X1 U420 ( .A(KEYINPUT109), .ZN(n431) );
  NOR2_X1 U421 ( .A1(n421), .A2(n420), .ZN(n419) );
  NOR2_X1 U422 ( .A1(n422), .A2(n494), .ZN(n421) );
  OR2_X1 U423 ( .A1(n440), .A2(n420), .ZN(n395) );
  XNOR2_X1 U424 ( .A(G107), .B(G104), .ZN(n452) );
  XNOR2_X1 U425 ( .A(KEYINPUT77), .B(G110), .ZN(n451) );
  XNOR2_X1 U426 ( .A(KEYINPUT16), .B(G122), .ZN(n482) );
  XOR2_X1 U427 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n458) );
  XNOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT80), .ZN(n457) );
  XNOR2_X1 U429 ( .A(KEYINPUT10), .B(G140), .ZN(n461) );
  AND2_X1 U430 ( .A1(n507), .A2(G221), .ZN(n443) );
  XNOR2_X1 U431 ( .A(G128), .B(G110), .ZN(n455) );
  OR2_X1 U432 ( .A1(n620), .A2(n390), .ZN(n384) );
  XNOR2_X1 U433 ( .A(n746), .B(n433), .ZN(n450) );
  XNOR2_X1 U434 ( .A(G146), .B(G140), .ZN(n433) );
  NAND2_X1 U435 ( .A1(n354), .A2(n373), .ZN(n607) );
  XNOR2_X1 U436 ( .A(n412), .B(n411), .ZN(n604) );
  XNOR2_X1 U437 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n411) );
  NAND2_X1 U438 ( .A1(n645), .A2(n492), .ZN(n397) );
  XNOR2_X1 U439 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U440 ( .A(n627), .B(n626), .ZN(n628) );
  INV_X1 U441 ( .A(KEYINPUT40), .ZN(n423) );
  NAND2_X1 U442 ( .A1(n534), .A2(n533), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n555), .B(KEYINPUT106), .ZN(n650) );
  NAND2_X1 U444 ( .A1(n554), .A2(n442), .ZN(n555) );
  XNOR2_X1 U445 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U446 ( .A(n645), .B(KEYINPUT62), .ZN(n646) );
  AND2_X1 U447 ( .A1(n439), .A2(n441), .ZN(n354) );
  AND2_X1 U448 ( .A1(n675), .A2(n685), .ZN(n355) );
  AND2_X1 U449 ( .A1(n402), .A2(n379), .ZN(n356) );
  NOR2_X1 U450 ( .A1(n583), .A2(n584), .ZN(n357) );
  INV_X1 U451 ( .A(KEYINPUT88), .ZN(n420) );
  XNOR2_X1 U452 ( .A(n607), .B(KEYINPUT38), .ZN(n672) );
  AND2_X1 U453 ( .A1(n750), .A2(n430), .ZN(n358) );
  NAND2_X1 U454 ( .A1(n437), .A2(n420), .ZN(n359) );
  XNOR2_X1 U455 ( .A(KEYINPUT73), .B(KEYINPUT39), .ZN(n360) );
  INV_X1 U456 ( .A(KEYINPUT74), .ZN(n409) );
  XNOR2_X1 U457 ( .A(n352), .B(n497), .ZN(n361) );
  XNOR2_X1 U458 ( .A(n595), .B(n497), .ZN(n605) );
  NAND2_X1 U459 ( .A1(n387), .A2(n383), .ZN(n362) );
  NAND2_X1 U460 ( .A1(n387), .A2(n383), .ZN(n363) );
  XNOR2_X1 U461 ( .A(n617), .B(KEYINPUT48), .ZN(n364) );
  BUF_X1 U462 ( .A(n610), .Z(n365) );
  NAND2_X1 U463 ( .A1(n387), .A2(n383), .ZN(n664) );
  XNOR2_X1 U464 ( .A(n617), .B(KEYINPUT48), .ZN(n751) );
  XNOR2_X1 U465 ( .A(n418), .B(KEYINPUT45), .ZN(n366) );
  XNOR2_X1 U466 ( .A(n418), .B(KEYINPUT45), .ZN(n727) );
  XNOR2_X1 U467 ( .A(n425), .B(KEYINPUT42), .ZN(n759) );
  NAND2_X1 U468 ( .A1(n667), .A2(n492), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n432), .B(n431), .ZN(n580) );
  XNOR2_X1 U470 ( .A(n473), .B(n398), .ZN(n645) );
  NAND2_X1 U471 ( .A1(n601), .A2(n689), .ZN(n412) );
  AND2_X2 U472 ( .A1(n378), .A2(n396), .ZN(n368) );
  NOR2_X1 U473 ( .A1(n596), .A2(n352), .ZN(n599) );
  NAND2_X1 U474 ( .A1(n509), .A2(KEYINPUT4), .ZN(n371) );
  NAND2_X1 U475 ( .A1(n369), .A2(n370), .ZN(n372) );
  NAND2_X1 U476 ( .A1(n371), .A2(n372), .ZN(n743) );
  INV_X1 U477 ( .A(n509), .ZN(n369) );
  AND2_X1 U478 ( .A1(n364), .A2(n358), .ZN(n377) );
  NOR2_X2 U479 ( .A1(n583), .A2(n400), .ZN(n399) );
  NAND2_X1 U480 ( .A1(n602), .A2(n560), .ZN(n432) );
  BUF_X1 U481 ( .A(n536), .Z(n559) );
  OR2_X1 U482 ( .A1(n625), .A2(n440), .ZN(n439) );
  AND2_X1 U483 ( .A1(n625), .A2(n494), .ZN(n374) );
  OR2_X1 U484 ( .A1(n625), .A2(n422), .ZN(n394) );
  INV_X1 U485 ( .A(n374), .ZN(n373) );
  NAND2_X1 U486 ( .A1(n381), .A2(n439), .ZN(n380) );
  NOR2_X1 U487 ( .A1(n374), .A2(n359), .ZN(n381) );
  AND2_X2 U488 ( .A1(n375), .A2(n388), .ZN(n387) );
  NAND2_X1 U489 ( .A1(n367), .A2(n427), .ZN(n375) );
  NAND2_X1 U490 ( .A1(n391), .A2(n389), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n377), .A2(n366), .ZN(n392) );
  AND2_X2 U492 ( .A1(n356), .A2(n616), .ZN(n617) );
  NOR2_X2 U493 ( .A1(n760), .A2(n759), .ZN(n615) );
  XNOR2_X2 U494 ( .A(n424), .B(n423), .ZN(n760) );
  NAND2_X1 U495 ( .A1(n394), .A2(n419), .ZN(n378) );
  INV_X1 U496 ( .A(n391), .ZN(n393) );
  NAND2_X1 U497 ( .A1(n427), .A2(n429), .ZN(n391) );
  NAND2_X1 U498 ( .A1(n393), .A2(n392), .ZN(n671) );
  NAND2_X1 U499 ( .A1(n386), .A2(n389), .ZN(n385) );
  INV_X1 U500 ( .A(n392), .ZN(n386) );
  NAND2_X1 U501 ( .A1(n605), .A2(n503), .ZN(n505) );
  OR2_X1 U502 ( .A1(n625), .A2(n395), .ZN(n396) );
  XNOR2_X2 U503 ( .A(n397), .B(G472), .ZN(n689) );
  XNOR2_X1 U504 ( .A(n479), .B(n480), .ZN(n398) );
  XNOR2_X1 U505 ( .A(n399), .B(n360), .ZN(n610) );
  NAND2_X1 U506 ( .A1(n401), .A2(n672), .ZN(n400) );
  INV_X1 U507 ( .A(n584), .ZN(n401) );
  NOR2_X1 U508 ( .A1(n406), .A2(n403), .ZN(n402) );
  NAND2_X1 U509 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U510 ( .A1(n643), .A2(KEYINPUT74), .ZN(n404) );
  NOR2_X1 U511 ( .A1(n410), .A2(n407), .ZN(n406) );
  NAND2_X1 U512 ( .A1(n408), .A2(n409), .ZN(n407) );
  XNOR2_X2 U513 ( .A(n415), .B(n454), .ZN(n602) );
  XNOR2_X2 U514 ( .A(n489), .B(n416), .ZN(n667) );
  INV_X1 U515 ( .A(n453), .ZN(n416) );
  XNOR2_X2 U516 ( .A(n489), .B(n417), .ZN(n625) );
  XNOR2_X2 U517 ( .A(n736), .B(n488), .ZN(n417) );
  XNOR2_X2 U518 ( .A(n472), .B(n734), .ZN(n489) );
  XNOR2_X2 U519 ( .A(n743), .B(G101), .ZN(n472) );
  NAND2_X1 U520 ( .A1(n636), .A2(n644), .ZN(n550) );
  NAND2_X1 U521 ( .A1(n544), .A2(n543), .ZN(n636) );
  NAND2_X1 U522 ( .A1(n494), .A2(n490), .ZN(n441) );
  INV_X1 U523 ( .A(n705), .ZN(n696) );
  NAND2_X1 U524 ( .A1(n610), .A2(n720), .ZN(n424) );
  NOR2_X1 U525 ( .A1(n705), .A2(n426), .ZN(n425) );
  INV_X1 U526 ( .A(n614), .ZN(n426) );
  NAND2_X1 U527 ( .A1(n727), .A2(n750), .ZN(n428) );
  OR2_X2 U528 ( .A1(n751), .A2(n430), .ZN(n429) );
  INV_X1 U529 ( .A(KEYINPUT2), .ZN(n430) );
  NOR2_X1 U530 ( .A1(n432), .A2(n689), .ZN(n561) );
  XNOR2_X2 U531 ( .A(n445), .B(n444), .ZN(n477) );
  XNOR2_X2 U532 ( .A(n434), .B(G143), .ZN(n509) );
  XNOR2_X2 U533 ( .A(G128), .B(KEYINPUT64), .ZN(n434) );
  NOR2_X1 U534 ( .A1(n438), .A2(n676), .ZN(n437) );
  INV_X1 U535 ( .A(n441), .ZN(n438) );
  AND2_X1 U536 ( .A1(n683), .A2(n686), .ZN(n442) );
  INV_X1 U537 ( .A(KEYINPUT92), .ZN(n446) );
  INV_X1 U538 ( .A(KEYINPUT81), .ZN(n447) );
  AND2_X1 U539 ( .A1(n720), .A2(n601), .ZN(n589) );
  XNOR2_X1 U540 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U541 ( .A(n450), .B(n449), .ZN(n453) );
  XNOR2_X1 U542 ( .A(n597), .B(KEYINPUT36), .ZN(n598) );
  INV_X1 U543 ( .A(KEYINPUT78), .ZN(n581) );
  XNOR2_X1 U544 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U545 ( .A(G134), .B(KEYINPUT70), .ZN(n444) );
  NAND2_X1 U546 ( .A1(G227), .A2(n755), .ZN(n448) );
  XNOR2_X1 U547 ( .A(n452), .B(n451), .ZN(n734) );
  INV_X1 U548 ( .A(G902), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT71), .B(G469), .Z(n454) );
  XNOR2_X1 U550 ( .A(n602), .B(KEYINPUT1), .ZN(n540) );
  XOR2_X1 U551 ( .A(G137), .B(G119), .Z(n456) );
  XNOR2_X1 U552 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U553 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U554 ( .A(n460), .B(n459), .Z(n463) );
  XNOR2_X2 U555 ( .A(G146), .B(G125), .ZN(n486) );
  XNOR2_X1 U556 ( .A(n744), .B(n443), .ZN(n462) );
  XNOR2_X1 U557 ( .A(n463), .B(n462), .ZN(n653) );
  NAND2_X1 U558 ( .A1(n653), .A2(n492), .ZN(n467) );
  XNOR2_X1 U559 ( .A(KEYINPUT15), .B(G902), .ZN(n619) );
  NAND2_X1 U560 ( .A1(n619), .A2(G234), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n464), .B(KEYINPUT20), .ZN(n468) );
  NAND2_X1 U562 ( .A1(n468), .A2(G217), .ZN(n465) );
  XNOR2_X1 U563 ( .A(KEYINPUT25), .B(n465), .ZN(n466) );
  XNOR2_X1 U564 ( .A(n467), .B(n466), .ZN(n585) );
  AND2_X1 U565 ( .A1(n468), .A2(G221), .ZN(n470) );
  XNOR2_X1 U566 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n469) );
  XNOR2_X1 U567 ( .A(n470), .B(n469), .ZN(n685) );
  INV_X1 U568 ( .A(n685), .ZN(n471) );
  OR2_X1 U569 ( .A1(n585), .A2(n471), .ZN(n682) );
  INV_X1 U570 ( .A(n682), .ZN(n560) );
  NAND2_X1 U571 ( .A1(n540), .A2(n560), .ZN(n556) );
  BUF_X1 U572 ( .A(n472), .Z(n473) );
  XOR2_X1 U573 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n475) );
  XNOR2_X1 U574 ( .A(G146), .B(KEYINPUT95), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U576 ( .A(n477), .B(n476), .Z(n480) );
  NAND2_X1 U577 ( .A1(n521), .A2(G210), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n483), .B(n478), .ZN(n479) );
  XNOR2_X1 U579 ( .A(n689), .B(KEYINPUT6), .ZN(n545) );
  XNOR2_X1 U580 ( .A(n481), .B(KEYINPUT33), .ZN(n704) );
  NAND2_X1 U581 ( .A1(n755), .A2(G224), .ZN(n484) );
  XNOR2_X1 U582 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U583 ( .A(n487), .B(n486), .ZN(n488) );
  INV_X1 U584 ( .A(n619), .ZN(n490) );
  NAND2_X1 U585 ( .A1(n492), .A2(n491), .ZN(n495) );
  NAND2_X1 U586 ( .A1(n495), .A2(G210), .ZN(n493) );
  XNOR2_X1 U587 ( .A(n493), .B(KEYINPUT90), .ZN(n494) );
  NAND2_X1 U588 ( .A1(n495), .A2(G214), .ZN(n611) );
  INV_X1 U589 ( .A(n611), .ZN(n676) );
  XNOR2_X1 U590 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n496) );
  XNOR2_X1 U591 ( .A(n496), .B(KEYINPUT67), .ZN(n497) );
  XOR2_X1 U592 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n499) );
  XNOR2_X1 U593 ( .A(n499), .B(n498), .ZN(n501) );
  NAND2_X1 U594 ( .A1(G952), .A2(n501), .ZN(n701) );
  NOR2_X1 U595 ( .A1(n701), .A2(G953), .ZN(n579) );
  NOR2_X1 U596 ( .A1(G898), .A2(n755), .ZN(n500) );
  XNOR2_X1 U597 ( .A(KEYINPUT91), .B(n500), .ZN(n738) );
  NAND2_X1 U598 ( .A1(G902), .A2(n501), .ZN(n576) );
  NOR2_X1 U599 ( .A1(n738), .A2(n576), .ZN(n502) );
  OR2_X1 U600 ( .A1(n579), .A2(n502), .ZN(n503) );
  XNOR2_X1 U601 ( .A(n505), .B(n504), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n704), .A2(n559), .ZN(n506) );
  XNOR2_X1 U603 ( .A(n506), .B(KEYINPUT34), .ZN(n534) );
  NAND2_X1 U604 ( .A1(n507), .A2(G217), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n509), .B(n508), .ZN(n516) );
  XNOR2_X1 U606 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U607 ( .A(n512), .B(KEYINPUT7), .Z(n514) );
  XNOR2_X1 U608 ( .A(G134), .B(G116), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n516), .B(n515), .ZN(n621) );
  NOR2_X1 U611 ( .A1(n621), .A2(G902), .ZN(n517) );
  XOR2_X1 U612 ( .A(n517), .B(G478), .Z(n565) );
  XNOR2_X1 U613 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U614 ( .A(n744), .B(n520), .Z(n529) );
  XOR2_X1 U615 ( .A(KEYINPUT97), .B(KEYINPUT99), .Z(n523) );
  NAND2_X1 U616 ( .A1(n521), .A2(G214), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n523), .B(n522), .ZN(n527) );
  XOR2_X1 U618 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n525) );
  XNOR2_X1 U619 ( .A(G122), .B(KEYINPUT12), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U621 ( .A(n527), .B(n526), .Z(n528) );
  XNOR2_X1 U622 ( .A(n529), .B(n528), .ZN(n657) );
  XNOR2_X1 U623 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n530) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n608) );
  XOR2_X1 U625 ( .A(KEYINPUT82), .B(n608), .Z(n533) );
  INV_X1 U626 ( .A(KEYINPUT35), .ZN(n535) );
  INV_X1 U627 ( .A(n536), .ZN(n538) );
  NOR2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n537) );
  XOR2_X1 U629 ( .A(KEYINPUT105), .B(n537), .Z(n675) );
  NAND2_X1 U630 ( .A1(n538), .A2(n355), .ZN(n539) );
  XNOR2_X1 U631 ( .A(n539), .B(KEYINPUT22), .ZN(n546) );
  BUF_X1 U632 ( .A(n546), .Z(n541) );
  INV_X1 U633 ( .A(n540), .ZN(n683) );
  INV_X1 U634 ( .A(n683), .ZN(n591) );
  NOR2_X1 U635 ( .A1(n541), .A2(n591), .ZN(n542) );
  XNOR2_X1 U636 ( .A(n542), .B(KEYINPUT108), .ZN(n544) );
  INV_X1 U637 ( .A(n585), .ZN(n686) );
  NOR2_X1 U638 ( .A1(n689), .A2(n686), .ZN(n543) );
  INV_X1 U639 ( .A(n545), .ZN(n588) );
  OR2_X2 U640 ( .A1(n546), .A2(n588), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n591), .A2(n585), .ZN(n547) );
  NOR2_X1 U642 ( .A1(n553), .A2(n547), .ZN(n549) );
  XOR2_X1 U643 ( .A(KEYINPUT83), .B(KEYINPUT32), .Z(n548) );
  XNOR2_X1 U644 ( .A(n549), .B(n548), .ZN(n642) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT44), .ZN(n574) );
  INV_X1 U646 ( .A(n556), .ZN(n557) );
  NAND2_X1 U647 ( .A1(n557), .A2(n689), .ZN(n692) );
  NOR2_X1 U648 ( .A1(n559), .A2(n692), .ZN(n558) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT31), .ZN(n639) );
  INV_X1 U650 ( .A(n559), .ZN(n562) );
  NAND2_X1 U651 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U652 ( .A(n563), .B(KEYINPUT96), .ZN(n712) );
  NAND2_X1 U653 ( .A1(n639), .A2(n712), .ZN(n570) );
  XOR2_X1 U654 ( .A(n564), .B(KEYINPUT101), .Z(n567) );
  INV_X1 U655 ( .A(n565), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n567), .A2(n568), .ZN(n566) );
  XNOR2_X2 U657 ( .A(n566), .B(KEYINPUT103), .ZN(n720) );
  NOR2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n716) );
  XOR2_X1 U659 ( .A(KEYINPUT104), .B(n569), .Z(n673) );
  NAND2_X1 U660 ( .A1(n570), .A2(n673), .ZN(n571) );
  NAND2_X1 U661 ( .A1(n650), .A2(n571), .ZN(n572) );
  XNOR2_X1 U662 ( .A(n572), .B(KEYINPUT107), .ZN(n573) );
  NAND2_X1 U663 ( .A1(n689), .A2(n611), .ZN(n575) );
  XNOR2_X1 U664 ( .A(KEYINPUT30), .B(n575), .ZN(n584) );
  OR2_X1 U665 ( .A1(n755), .A2(n576), .ZN(n577) );
  NOR2_X1 U666 ( .A1(G900), .A2(n577), .ZN(n578) );
  NOR2_X1 U667 ( .A1(n579), .A2(n578), .ZN(n587) );
  NOR2_X2 U668 ( .A1(n580), .A2(n587), .ZN(n582) );
  XNOR2_X1 U669 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U670 ( .A1(n365), .A2(n716), .ZN(n726) );
  NAND2_X1 U671 ( .A1(n685), .A2(n585), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n589), .A2(n588), .ZN(n596) );
  OR2_X1 U673 ( .A1(n596), .A2(n676), .ZN(n590) );
  NOR2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U675 ( .A(n592), .B(KEYINPUT43), .ZN(n594) );
  INV_X1 U676 ( .A(n607), .ZN(n593) );
  OR2_X1 U677 ( .A1(n594), .A2(n593), .ZN(n633) );
  AND2_X1 U678 ( .A1(n726), .A2(n633), .ZN(n750) );
  XNOR2_X1 U679 ( .A(KEYINPUT87), .B(KEYINPUT112), .ZN(n597) );
  NOR2_X1 U680 ( .A1(n683), .A2(n600), .ZN(n724) );
  INV_X1 U681 ( .A(n602), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n614) );
  AND2_X1 U683 ( .A1(n361), .A2(n614), .ZN(n721) );
  NAND2_X1 U684 ( .A1(n673), .A2(n721), .ZN(n606) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U686 ( .A1(n357), .A2(n609), .ZN(n643) );
  XOR2_X1 U687 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n613) );
  AND2_X1 U688 ( .A1(n675), .A2(n672), .ZN(n679) );
  NAND2_X1 U689 ( .A1(n679), .A2(n611), .ZN(n612) );
  XOR2_X1 U690 ( .A(n613), .B(n612), .Z(n705) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT46), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n430), .A2(KEYINPUT84), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n620) );
  INV_X1 U694 ( .A(n621), .ZN(n622) );
  INV_X1 U695 ( .A(G952), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n623), .A2(G953), .ZN(n660) );
  INV_X1 U697 ( .A(KEYINPUT120), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n363), .A2(G210), .ZN(n629) );
  BUF_X1 U699 ( .A(n625), .Z(n627) );
  XNOR2_X1 U700 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n630), .A2(n660), .ZN(n632) );
  INV_X1 U703 ( .A(KEYINPUT56), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n632), .B(n631), .ZN(G51) );
  XNOR2_X1 U705 ( .A(n633), .B(G140), .ZN(G42) );
  INV_X1 U706 ( .A(n712), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n634), .A2(n720), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n635), .B(G104), .ZN(G6) );
  XNOR2_X1 U709 ( .A(n636), .B(G110), .ZN(G12) );
  INV_X1 U710 ( .A(n639), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n637), .A2(n720), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n638), .B(G113), .ZN(G15) );
  INV_X1 U713 ( .A(n716), .ZN(n711) );
  NOR2_X1 U714 ( .A1(n639), .A2(n711), .ZN(n640) );
  XOR2_X1 U715 ( .A(G116), .B(n640), .Z(G18) );
  XNOR2_X1 U716 ( .A(G119), .B(KEYINPUT127), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(G21) );
  XOR2_X1 U718 ( .A(G143), .B(n643), .Z(G45) );
  XNOR2_X1 U719 ( .A(n644), .B(G122), .ZN(G24) );
  NAND2_X1 U720 ( .A1(n664), .A2(G472), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n648), .A2(n660), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(KEYINPUT63), .ZN(G57) );
  BUF_X1 U724 ( .A(n650), .Z(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(G101), .ZN(G3) );
  NAND2_X1 U726 ( .A1(n363), .A2(G217), .ZN(n652) );
  XOR2_X1 U727 ( .A(n653), .B(n652), .Z(n654) );
  NOR2_X1 U728 ( .A1(n654), .A2(n341), .ZN(G66) );
  NAND2_X1 U729 ( .A1(n664), .A2(G475), .ZN(n659) );
  XNOR2_X1 U730 ( .A(KEYINPUT66), .B(KEYINPUT119), .ZN(n655) );
  XOR2_X1 U731 ( .A(n655), .B(KEYINPUT59), .Z(n656) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n663) );
  XOR2_X1 U734 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n362), .A2(G469), .ZN(n669) );
  XNOR2_X1 U737 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(KEYINPUT58), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n670), .A2(n341), .ZN(G54) );
  AND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n704), .A2(n680), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(KEYINPUT115), .ZN(n698) );
  NAND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT50), .ZN(n691) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U751 ( .A(KEYINPUT49), .B(n687), .Z(n688) );
  NOR2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n694), .Z(n695) );
  NAND2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U758 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n699) );
  XNOR2_X1 U759 ( .A(n700), .B(n699), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U761 ( .A1(n703), .A2(G953), .ZN(n707) );
  OR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U763 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U764 ( .A1(n671), .A2(n708), .ZN(n710) );
  XOR2_X1 U765 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n709) );
  XNOR2_X1 U766 ( .A(n710), .B(n709), .ZN(G75) );
  XOR2_X1 U767 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n714) );
  NOR2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U769 ( .A(n714), .B(n713), .Z(n715) );
  XNOR2_X1 U770 ( .A(G107), .B(n715), .ZN(G9) );
  XOR2_X1 U771 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n718) );
  NAND2_X1 U772 ( .A1(n721), .A2(n716), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U774 ( .A(G128), .B(n719), .Z(G30) );
  NAND2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U776 ( .A(n722), .B(KEYINPUT114), .ZN(n723) );
  XNOR2_X1 U777 ( .A(G146), .B(n723), .ZN(G48) );
  XNOR2_X1 U778 ( .A(G125), .B(n724), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n725), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U780 ( .A(G134), .B(n726), .ZN(G36) );
  AND2_X1 U781 ( .A1(n366), .A2(n755), .ZN(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n729) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U785 ( .A1(G898), .A2(n730), .ZN(n731) );
  XOR2_X1 U786 ( .A(KEYINPUT122), .B(n731), .Z(n732) );
  NOR2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n742) );
  XNOR2_X1 U788 ( .A(n734), .B(KEYINPUT123), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(G101), .B(n737), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n740), .B(KEYINPUT124), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n353), .B(n744), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(n752) );
  XOR2_X1 U796 ( .A(G227), .B(n752), .Z(n747) );
  NAND2_X1 U797 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U798 ( .A1(G953), .A2(n748), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n749), .B(KEYINPUT126), .ZN(n758) );
  NAND2_X1 U800 ( .A1(n364), .A2(n750), .ZN(n754) );
  XNOR2_X1 U801 ( .A(KEYINPUT125), .B(n752), .ZN(n753) );
  XNOR2_X1 U802 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U805 ( .A(G137), .B(n759), .Z(G39) );
  XOR2_X1 U806 ( .A(n760), .B(G131), .Z(G33) );
endmodule

