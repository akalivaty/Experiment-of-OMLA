//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(new_n470), .B1(G113), .B2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .A3(G125), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n465), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(new_n479), .A3(new_n464), .A4(new_n468), .ZN(new_n480));
  INV_X1    g055(.A(G137), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n474), .A2(new_n482), .ZN(G160));
  INV_X1    g058(.A(new_n480), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT70), .Z(new_n488));
  NAND4_X1  g063(.A1(new_n478), .A2(new_n479), .A3(G2105), .A4(new_n468), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n485), .B(new_n488), .C1(G124), .C2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n478), .A2(new_n479), .A3(new_n493), .A4(new_n468), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n472), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n464), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n489), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n496), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT71), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(new_n502), .A3(KEYINPUT5), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(G62), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(KEYINPUT72), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n508), .A2(new_n517), .A3(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n514), .B1(new_n519), .B2(G651), .ZN(G166));
  INV_X1    g095(.A(new_n510), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n513), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT73), .B(G51), .Z(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n523), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n510), .A2(new_n535), .B1(new_n536), .B2(new_n513), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n533), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n510), .A2(new_n541), .B1(new_n542), .B2(new_n513), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n505), .A2(new_n507), .ZN(new_n557));
  INV_X1    g132(.A(new_n503), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n557), .A2(G91), .A3(new_n558), .A4(new_n509), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT77), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n508), .A2(new_n561), .A3(G91), .A4(new_n509), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(G65), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  INV_X1    g141(.A(new_n564), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n508), .B2(G65), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n560), .B(new_n562), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n513), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n509), .A2(new_n574), .A3(G53), .A4(G543), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n572), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n560), .A2(new_n562), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n533), .B1(new_n568), .B2(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n563), .A2(new_n564), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n572), .A2(new_n575), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n580), .A2(new_n593), .ZN(G299));
  INV_X1    g169(.A(G171), .ZN(G301));
  INV_X1    g170(.A(G166), .ZN(G303));
  NAND3_X1  g171(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n521), .A2(G87), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G288));
  AND2_X1   g176(.A1(KEYINPUT6), .A2(G651), .ZN(new_n602));
  NOR2_X1   g177(.A1(KEYINPUT6), .A2(G651), .ZN(new_n603));
  OAI211_X1 g178(.A(G48), .B(G543), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT82), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n509), .A2(new_n606), .A3(G48), .A4(G543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n533), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n557), .A2(G86), .A3(new_n558), .A4(new_n509), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT81), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n508), .A2(new_n613), .A3(G86), .A4(new_n509), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(G305));
  INV_X1    g192(.A(G85), .ZN(new_n618));
  INV_X1    g193(.A(G47), .ZN(new_n619));
  OAI22_X1  g194(.A1(new_n510), .A2(new_n618), .B1(new_n619), .B2(new_n513), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(new_n533), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n620), .B1(new_n622), .B2(KEYINPUT83), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(KEYINPUT83), .B2(new_n622), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n521), .A2(G92), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n508), .A2(G66), .ZN(new_n629));
  INV_X1    g204(.A(G79), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n502), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n631), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n625), .B1(new_n633), .B2(G868), .ZN(G284));
  OAI21_X1  g209(.A(new_n625), .B1(new_n633), .B2(G868), .ZN(G321));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(G299), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(G168), .ZN(G297));
  OAI21_X1  g213(.A(new_n637), .B1(new_n636), .B2(G168), .ZN(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n633), .B1(new_n640), .B2(G860), .ZN(G148));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n633), .A2(new_n640), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(G868), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n550), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n642), .A3(G868), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(G323));
  XOR2_X1   g222(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n648));
  XNOR2_X1  g223(.A(G323), .B(new_n648), .ZN(G282));
  INV_X1    g224(.A(G135), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n480), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  INV_X1    g228(.A(G111), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(G2105), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n490), .B2(G123), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT88), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(G2096), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(G2096), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n472), .A2(new_n475), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT13), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G2100), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2435), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT90), .B(G2438), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2427), .B(G2430), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(KEYINPUT14), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2443), .B(G2446), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2451), .B(G2454), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(G14), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n681), .B2(new_n678), .ZN(G401));
  XOR2_X1   g258(.A(G2067), .B(G2678), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT18), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(KEYINPUT17), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n691), .B(new_n688), .C1(new_n685), .C2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n685), .A3(new_n687), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G2096), .B(G2100), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  XOR2_X1   g278(.A(G1961), .B(G1966), .Z(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT20), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n702), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n702), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT92), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(G1986), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n714), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n714), .B2(new_n718), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n699), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n721), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n723), .A2(new_n719), .A3(new_n698), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(G229));
  NAND2_X1  g300(.A1(new_n484), .A2(G140), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n490), .A2(G128), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n464), .A2(G116), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT95), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G105), .B2(new_n475), .ZN(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n489), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G141), .B2(new_n484), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n733), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT27), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G1996), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(G1996), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n738), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G21), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G168), .B2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n758));
  OR2_X1    g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n757), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n755), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(G29), .A2(G33), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n484), .A2(G139), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  AOI22_X1  g341(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n766), .C1(new_n464), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(new_n733), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n442), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n754), .A2(G1966), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n762), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT24), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT24), .ZN(new_n775));
  AOI22_X1  g350(.A1(G160), .A2(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G2084), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  INV_X1    g353(.A(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n779), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n777), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n733), .A2(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n733), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(new_n443), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n781), .A2(G1961), .B1(new_n776), .B2(G2084), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n772), .A2(new_n783), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n628), .A2(new_n632), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n779), .ZN(new_n790));
  INV_X1    g365(.A(G1348), .ZN(new_n791));
  NOR2_X1   g366(.A1(G4), .A2(G16), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n769), .A2(new_n442), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n658), .A2(G29), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n793), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n752), .A2(new_n788), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(G162), .A2(G29), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G29), .B2(G35), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2090), .ZN(new_n804));
  NAND2_X1  g379(.A1(G299), .A2(G16), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n779), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n779), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n550), .B2(new_n779), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1341), .Z(new_n813));
  NAND4_X1  g388(.A1(new_n799), .A2(new_n804), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n779), .A2(G23), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n779), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT33), .B(G1976), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(G166), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G16), .B2(G22), .ZN(new_n823));
  INV_X1    g398(.A(G1971), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n779), .A2(G6), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n616), .B2(new_n779), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT32), .B(G1981), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n818), .B2(new_n820), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n827), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n827), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n733), .A2(G25), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n484), .A2(G131), .ZN(new_n837));
  INV_X1    g412(.A(G119), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n464), .A2(G107), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n489), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n836), .B1(new_n842), .B2(new_n733), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT35), .B(G1991), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n843), .B(new_n844), .Z(new_n845));
  INV_X1    g420(.A(G1986), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n779), .A2(G24), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G290), .B2(G16), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n845), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n846), .B2(new_n848), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n834), .A2(new_n835), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n834), .A2(new_n853), .A3(new_n835), .A4(new_n850), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n814), .B1(new_n852), .B2(new_n854), .ZN(G311));
  NOR2_X1   g430(.A1(G311), .A2(KEYINPUT98), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n857));
  AOI211_X1 g432(.A(new_n857), .B(new_n814), .C1(new_n852), .C2(new_n854), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(G150));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  INV_X1    g435(.A(G55), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n510), .A2(new_n860), .B1(new_n861), .B2(new_n513), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT100), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n533), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n789), .A2(new_n640), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n549), .A2(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n863), .A2(new_n544), .A3(new_n865), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n872), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n869), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(KEYINPUT101), .A3(new_n877), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n868), .B1(new_n885), .B2(new_n886), .ZN(G145));
  XNOR2_X1  g462(.A(new_n658), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G162), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n768), .A2(KEYINPUT104), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n747), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n730), .ZN(new_n892));
  INV_X1    g467(.A(new_n500), .ZN(new_n893));
  AOI221_X4 g468(.A(KEYINPUT103), .B1(new_n472), .B2(new_n495), .C1(new_n494), .C2(KEYINPUT4), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n472), .A2(new_n495), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n893), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n892), .B(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n842), .B(new_n664), .Z(new_n902));
  INV_X1    g477(.A(G130), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n464), .A2(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n489), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(G142), .B2(new_n484), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n902), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n889), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n901), .A2(new_n908), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n901), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n901), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n889), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g493(.A(new_n875), .B(new_n643), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n789), .B1(new_n580), .B2(new_n593), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n591), .A2(new_n592), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n633), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT41), .B1(new_n920), .B2(new_n923), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n925), .B1(new_n929), .B2(new_n919), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G290), .B(new_n616), .ZN(new_n933));
  XNOR2_X1  g508(.A(G166), .B(new_n816), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n925), .B(KEYINPUT107), .C1(new_n919), .C2(new_n929), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n866), .A2(new_n636), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(G331));
  XNOR2_X1  g519(.A(G171), .B(G286), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n873), .A2(new_n874), .A3(new_n946), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n546), .A2(new_n548), .B1(new_n863), .B2(new_n865), .ZN(new_n948));
  INV_X1    g523(.A(new_n874), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT41), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n924), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n951), .B1(new_n953), .B2(new_n926), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n924), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n935), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n951), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n927), .B2(new_n928), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n933), .B(new_n934), .Z(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n955), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n957), .A2(new_n961), .A3(new_n966), .A4(new_n962), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(KEYINPUT44), .A3(new_n967), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(KEYINPUT118), .ZN(new_n974));
  INV_X1    g549(.A(G1976), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(G288), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G40), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n474), .A2(new_n977), .A3(new_n482), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n899), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT114), .B(G8), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n598), .A2(new_n599), .A3(G1976), .A4(new_n600), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n976), .A2(new_n980), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT52), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n896), .A2(new_n897), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT103), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n496), .A2(new_n895), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n990), .B2(new_n893), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n991), .B2(new_n978), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n610), .A2(new_n615), .A3(G1981), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n506), .B1(KEYINPUT5), .B2(new_n502), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n504), .A2(KEYINPUT71), .A3(G543), .ZN(new_n997));
  OAI211_X1 g572(.A(G61), .B(new_n558), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G73), .A2(G543), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n1000), .A2(G651), .B1(new_n605), .B2(new_n607), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n712), .B1(new_n1001), .B2(new_n611), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1001), .A2(new_n712), .A3(new_n612), .A4(new_n614), .ZN(new_n1005));
  INV_X1    g580(.A(new_n611), .ZN(new_n1006));
  OAI21_X1  g581(.A(G1981), .B1(new_n610), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT115), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n994), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n984), .B(new_n986), .C1(new_n1004), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(G166), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n533), .B1(new_n516), .B2(new_n518), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT55), .B(G8), .C1(new_n1015), .C2(new_n514), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n979), .B1(new_n496), .B2(new_n500), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n978), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n991), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n899), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n978), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1023), .A2(new_n1024), .B1(new_n1028), .B2(new_n824), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1018), .B1(new_n1029), .B2(new_n1013), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n899), .B2(new_n979), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n978), .B1(new_n1026), .B2(new_n1019), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n469), .A2(new_n470), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G113), .A2(G2104), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n473), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G2105), .ZN(new_n1038));
  INV_X1    g613(.A(new_n482), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(G40), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(KEYINPUT50), .B2(new_n1019), .ZN(new_n1041));
  INV_X1    g616(.A(G2084), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n899), .A2(new_n1022), .A3(new_n979), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI211_X1 g619(.A(G286), .B(new_n981), .C1(new_n1034), .C2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1011), .A2(new_n1030), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT63), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G288), .A2(G1976), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n980), .A2(new_n982), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n994), .B2(new_n1008), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1008), .A2(new_n994), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1054), .B2(new_n995), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1049), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT116), .A3(new_n1005), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n992), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1047), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1019), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1040), .B1(new_n1061), .B2(new_n1022), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1062), .B(new_n1063), .C1(new_n991), .C2(new_n1022), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1022), .B1(new_n899), .B2(new_n979), .ZN(new_n1065));
  OAI211_X1 g640(.A(G160), .B(G40), .C1(KEYINPUT50), .C2(new_n1019), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT117), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1067), .A3(new_n1024), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1028), .A2(new_n824), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n981), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1060), .B(new_n1045), .C1(new_n1070), .C2(new_n1017), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1069), .B1(G2090), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1014), .A2(new_n1074), .A3(new_n1016), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1073), .A2(new_n1076), .A3(G8), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1010), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n974), .B1(new_n1059), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1017), .B1(new_n1081), .B2(new_n982), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1045), .A2(new_n1060), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1011), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(KEYINPUT118), .A3(new_n1058), .A4(new_n1047), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n899), .A2(new_n979), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n1040), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1072), .A2(new_n791), .B1(new_n1089), .B2(new_n737), .ZN(new_n1090));
  OR3_X1    g665(.A1(new_n1090), .A2(KEYINPUT120), .A3(new_n789), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n809), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1025), .A2(new_n978), .A3(new_n1027), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n586), .B2(new_n590), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n587), .A2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n570), .A2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1097), .A2(new_n1099), .A3(KEYINPUT119), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT57), .B1(new_n570), .B2(new_n578), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n572), .B2(new_n575), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n586), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1095), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT120), .B1(new_n1090), .B2(new_n789), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1091), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1102), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1090), .A2(KEYINPUT60), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n899), .A2(new_n1022), .A3(new_n979), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n791), .B1(new_n1114), .B2(new_n1021), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n991), .A2(new_n737), .A3(new_n978), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n633), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1117), .B2(new_n633), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n789), .A4(new_n1116), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1113), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n549), .B1(new_n1126), .B2(KEYINPUT59), .ZN(new_n1127));
  INV_X1    g702(.A(G1996), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1025), .A2(new_n1128), .A3(new_n978), .A4(new_n1027), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n980), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1126), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g712(.A(new_n1127), .B1(new_n1126), .B2(KEYINPUT59), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1106), .A2(new_n1139), .A3(new_n1111), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1137), .B(new_n1138), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1112), .B1(new_n1125), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1081), .A2(new_n982), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1018), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1029), .A2(new_n1013), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1014), .A2(new_n1074), .A3(new_n1016), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(new_n1075), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1010), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1034), .A2(new_n1044), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(G286), .A3(new_n982), .ZN(new_n1151));
  NOR2_X1   g726(.A1(G168), .A2(new_n981), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1013), .B1(new_n1034), .B2(new_n1044), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1151), .B(KEYINPUT51), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n982), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1152), .A2(KEYINPUT51), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1145), .A2(new_n1149), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1028), .B2(G2078), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1072), .A2(new_n778), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1163));
  OR3_X1    g738(.A1(new_n1032), .A2(new_n1033), .A3(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(G171), .B(KEYINPUT54), .Z(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1032), .A2(new_n1163), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1167), .A2(new_n978), .A3(new_n1025), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1160), .A2(new_n1168), .A3(new_n1161), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1165), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT125), .B1(new_n1158), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1078), .A2(new_n1011), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(new_n1082), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1172), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1143), .A2(new_n1174), .A3(new_n1179), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1177), .A2(KEYINPUT62), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(KEYINPUT62), .ZN(new_n1182));
  AOI21_X1  g757(.A(G301), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1176), .A4(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1087), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G290), .A2(G1986), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT109), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1032), .A2(new_n978), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(G1986), .A3(G290), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT110), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n730), .B(G2067), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT112), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1195), .B1(new_n1128), .B2(new_n747), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1189), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1189), .A2(KEYINPUT111), .A3(new_n1128), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT111), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n1188), .B2(G1996), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n747), .ZN(new_n1202));
  INV_X1    g777(.A(new_n842), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1203), .A2(new_n844), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1203), .A2(new_n844), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1189), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1197), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1193), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1185), .A2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1201), .A2(KEYINPUT46), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT127), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT47), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1188), .B1(new_n1195), .B2(new_n747), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1201), .B2(KEYINPUT46), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1212), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1190), .B(KEYINPUT48), .Z(new_n1217));
  OAI22_X1  g792(.A1(new_n1215), .A2(new_n1216), .B1(new_n1217), .B2(new_n1207), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1197), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1219));
  OR2_X1    g794(.A1(new_n730), .A2(G2067), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1188), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT126), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1209), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g799(.A1(G401), .A2(G227), .A3(new_n462), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n722), .A2(new_n724), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n911), .B2(new_n916), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n1228), .A2(new_n968), .A3(new_n970), .ZN(G225));
  INV_X1    g803(.A(G225), .ZN(G308));
endmodule


