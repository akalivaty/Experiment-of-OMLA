//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(G237), .A2(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G143), .A3(G214), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n187), .B1(new_n195), .B2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  AOI211_X1 g011(.A(KEYINPUT86), .B(new_n197), .C1(new_n192), .C2(new_n194), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT17), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n202), .B1(new_n206), .B2(new_n200), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(G146), .B(new_n202), .C1(new_n206), .C2(new_n200), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AND4_X1   g026(.A1(G143), .A2(new_n188), .A3(new_n189), .A4(G214), .ZN(new_n213));
  AOI21_X1  g027(.A(G143), .B1(new_n193), .B2(G214), .ZN(new_n214));
  OAI21_X1  g028(.A(G131), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT86), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n195), .A2(new_n187), .A3(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n192), .A2(new_n197), .A3(new_n194), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT85), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n192), .A2(KEYINPUT85), .A3(new_n197), .A4(new_n194), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n216), .A2(new_n217), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n199), .B(new_n212), .C1(new_n222), .C2(KEYINPUT17), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT18), .A2(G131), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n195), .B(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT75), .B1(new_n206), .B2(G146), .ZN(new_n227));
  XNOR2_X1  g041(.A(G125), .B(G140), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n208), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n227), .A2(new_n230), .B1(G146), .B2(new_n206), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G113), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(G104), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n236), .B(KEYINPUT88), .Z(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n223), .A2(new_n233), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n236), .B1(new_n240), .B2(KEYINPUT89), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n220), .A2(new_n221), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n196), .A2(new_n198), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n216), .A2(new_n217), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n211), .B1(new_n246), .B2(KEYINPUT17), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n232), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n239), .B1(new_n241), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(G475), .B1(new_n251), .B2(G902), .ZN(new_n252));
  INV_X1    g066(.A(new_n236), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT19), .B1(new_n228), .B2(KEYINPUT87), .ZN(new_n254));
  AND4_X1   g068(.A1(KEYINPUT87), .A2(new_n203), .A3(new_n205), .A4(KEYINPUT19), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n208), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n210), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n242), .B2(new_n243), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n253), .B1(new_n258), .B2(new_n232), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n238), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G475), .A2(G902), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n260), .A2(new_n266), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n189), .A2(G952), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(G234), .B2(G237), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n271), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT21), .B(G898), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT9), .B(G234), .ZN(new_n276));
  INV_X1    g090(.A(G217), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(G953), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT90), .ZN(new_n280));
  INV_X1    g094(.A(G122), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G122), .ZN(new_n284));
  INV_X1    g098(.A(G107), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n282), .B2(new_n284), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n283), .A2(G122), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n281), .A2(G116), .ZN(new_n290));
  OAI21_X1  g104(.A(G107), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT90), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n191), .A2(G128), .ZN(new_n294));
  OAI21_X1  g108(.A(G134), .B1(new_n294), .B2(KEYINPUT13), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n191), .A2(G128), .ZN(new_n296));
  INV_X1    g110(.A(G128), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT13), .A4(G134), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n288), .A2(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT14), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n283), .A3(G122), .ZN(new_n304));
  OAI21_X1  g118(.A(G107), .B1(new_n304), .B2(KEYINPUT91), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT14), .B1(new_n281), .B2(G116), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n281), .A2(KEYINPUT14), .A3(G116), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT91), .B1(new_n283), .B2(G122), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G134), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n299), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n296), .A2(new_n298), .A3(G134), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n292), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n279), .B1(new_n302), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n300), .A2(new_n301), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n286), .A2(new_n287), .A3(new_n280), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT90), .B1(new_n291), .B2(new_n292), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n306), .A2(new_n304), .A3(KEYINPUT91), .A4(new_n282), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n321), .B(G107), .C1(KEYINPUT91), .C2(new_n304), .ZN(new_n322));
  AOI21_X1  g136(.A(G134), .B1(new_n296), .B2(new_n298), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n286), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n313), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n325), .A3(new_n278), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT92), .B(new_n279), .C1(new_n302), .C2(new_n315), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n328), .A2(KEYINPUT93), .A3(new_n271), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G478), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n331), .A2(KEYINPUT15), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n252), .A2(new_n268), .A3(new_n275), .A4(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G221), .ZN(new_n335));
  INV_X1    g149(.A(new_n276), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n271), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT64), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n208), .A3(G143), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n191), .A2(G146), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n191), .A2(G146), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n345));
  OAI21_X1  g159(.A(G128), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n297), .A2(KEYINPUT1), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n339), .A2(new_n341), .A3(new_n342), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n235), .B2(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n285), .A2(KEYINPUT3), .A3(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G101), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n285), .B2(G104), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n235), .A2(KEYINPUT79), .A3(G107), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT80), .B1(new_n285), .B2(G104), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n285), .A2(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n285), .A2(KEYINPUT80), .A3(G104), .ZN(new_n363));
  OAI21_X1  g177(.A(G101), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n359), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n345), .B1(G143), .B2(new_n208), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n208), .A2(G143), .ZN(new_n368));
  OAI22_X1  g182(.A1(new_n367), .A2(new_n297), .B1(new_n344), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n369), .A2(new_n349), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT66), .ZN(new_n373));
  INV_X1    g187(.A(G137), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G134), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(G134), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n373), .A2(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n311), .A2(G137), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT67), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT66), .B1(new_n374), .B2(G134), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n378), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n377), .B1(new_n311), .B2(G137), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n373), .A2(new_n311), .A3(G137), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n376), .B1(new_n389), .B2(new_n377), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT67), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(G131), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT68), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n388), .A2(new_n390), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n197), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n385), .A2(new_n391), .A3(new_n393), .A4(G131), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n372), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n372), .A2(KEYINPUT12), .A3(new_n396), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G140), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n189), .A2(G227), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n285), .A2(KEYINPUT3), .A3(G104), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT3), .B1(new_n285), .B2(G104), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n357), .B(new_n358), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G101), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT0), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n297), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n297), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(new_n414), .C1(new_n344), .C2(new_n368), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n408), .A2(new_n418), .A3(G101), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n410), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n347), .A2(new_n349), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n366), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n364), .A2(new_n359), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n369), .B2(new_n349), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n420), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n396), .A2(new_n397), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n405), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n402), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n396), .A2(new_n397), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n423), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n365), .A2(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n434), .A3(new_n420), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n405), .ZN(new_n437));
  AOI211_X1 g251(.A(G469), .B(G902), .C1(new_n430), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n405), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n400), .A2(new_n401), .B1(new_n427), .B2(new_n428), .ZN(new_n441));
  OAI211_X1 g255(.A(G469), .B(new_n440), .C1(new_n441), .C2(new_n439), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n271), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n338), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(G119), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n283), .A2(G119), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT2), .B(G113), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n453), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT70), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT70), .ZN(new_n458));
  INV_X1    g272(.A(new_n456), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n410), .A2(new_n457), .A3(new_n460), .A4(new_n419), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g276(.A(G113), .B1(new_n450), .B2(KEYINPUT5), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n454), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n424), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G122), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n461), .A2(new_n466), .A3(new_n468), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n369), .A2(new_n349), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G125), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n204), .B1(new_n415), .B2(new_n416), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G224), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G953), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n476), .B(new_n478), .Z(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n467), .A2(new_n480), .A3(new_n469), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n424), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n465), .B1(new_n366), .B2(KEYINPUT81), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n468), .B(KEYINPUT8), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT7), .B1(new_n477), .B2(G953), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n474), .B2(new_n475), .ZN(new_n490));
  OR3_X1    g304(.A1(new_n474), .A2(new_n475), .A3(new_n489), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n492), .B2(new_n471), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n482), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n482), .B2(new_n493), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n448), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT83), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(new_n448), .C1(new_n497), .C2(new_n498), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n334), .B(new_n447), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n277), .B1(G234), .B2(new_n271), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT74), .B1(new_n449), .B2(G128), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT74), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n297), .A3(G119), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n449), .A2(G128), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT24), .B(G110), .Z(new_n511));
  NAND3_X1  g325(.A1(new_n297), .A2(KEYINPUT23), .A3(G119), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n449), .A2(G128), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n509), .B(new_n512), .C1(new_n513), .C2(KEYINPUT23), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n510), .A2(new_n511), .B1(new_n514), .B2(G110), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n227), .A2(new_n230), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n210), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(new_n519), .A3(new_n516), .A4(new_n210), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n510), .A2(new_n511), .B1(new_n514), .B2(G110), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n211), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT22), .B(G137), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n527), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT77), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n505), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n528), .A2(new_n537), .A3(new_n530), .A4(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n528), .A2(new_n530), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n504), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT78), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OR3_X1    g357(.A1(new_n540), .A2(KEYINPUT78), .A3(new_n542), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n396), .A2(new_n417), .A3(new_n397), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n378), .A2(new_n382), .A3(new_n197), .A4(new_n384), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n379), .B2(new_n375), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n473), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n547), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n457), .A2(new_n460), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n396), .A2(new_n417), .A3(new_n397), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT30), .A3(new_n551), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n555), .A3(new_n551), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n193), .A2(G210), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(KEYINPUT27), .Z(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT26), .B(G101), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n562), .B(new_n563), .Z(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n559), .A2(KEYINPUT71), .A3(new_n560), .A4(new_n564), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT31), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n570));
  AND4_X1   g384(.A1(new_n559), .A2(new_n560), .A3(new_n564), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n551), .B(KEYINPUT69), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n555), .B1(new_n572), .B2(new_n557), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n557), .A2(new_n575), .A3(new_n555), .A4(new_n551), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n573), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n564), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n569), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n581), .A2(G472), .A3(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n555), .B1(new_n557), .B2(new_n551), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n574), .B2(new_n576), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n564), .A2(KEYINPUT29), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n559), .A2(new_n560), .ZN(new_n590));
  INV_X1    g404(.A(new_n564), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT73), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n593), .B(new_n564), .C1(new_n559), .C2(new_n560), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT29), .B1(new_n577), .B2(new_n564), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n589), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G472), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n583), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(G472), .A2(G902), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT32), .B1(new_n580), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n503), .B(new_n546), .C1(new_n599), .C2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND2_X1  g417(.A1(new_n580), .A2(new_n600), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n447), .A2(new_n545), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n569), .B2(new_n579), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n604), .B(new_n605), .C1(new_n598), .C2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n328), .A2(new_n608), .A3(new_n329), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n316), .A2(new_n326), .A3(KEYINPUT33), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n331), .A2(G902), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n328), .A2(new_n271), .A3(new_n329), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n331), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT94), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n252), .A2(new_n268), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n482), .A2(new_n493), .A3(new_n495), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n495), .B1(new_n482), .B2(new_n493), .ZN(new_n623));
  INV_X1    g437(.A(new_n448), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n274), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n607), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NAND2_X1  g443(.A1(new_n580), .A2(new_n271), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(G472), .B1(new_n600), .B2(new_n580), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT95), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n260), .A2(new_n263), .A3(new_n261), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n265), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n333), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n263), .B1(new_n260), .B2(new_n261), .ZN(new_n636));
  INV_X1    g450(.A(new_n261), .ZN(new_n637));
  AOI211_X1 g451(.A(new_n264), .B(new_n637), .C1(new_n238), .C2(new_n259), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT95), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n252), .A2(new_n634), .A3(new_n635), .A4(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n625), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n631), .A2(new_n605), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT96), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR3_X1   g459(.A1(new_n524), .A2(KEYINPUT36), .A3(new_n527), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n527), .A2(KEYINPUT36), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n521), .B2(new_n523), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n541), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n649), .A2(KEYINPUT97), .A3(new_n541), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n539), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n631), .A2(new_n503), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AND3_X1   g473(.A1(new_n652), .A2(new_n539), .A3(new_n653), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n482), .A2(new_n493), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n494), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n448), .A3(new_n621), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n442), .A2(new_n445), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n430), .A2(new_n437), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n443), .A3(new_n271), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n337), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n270), .B1(new_n272), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT100), .Z(new_n671));
  AND4_X1   g485(.A1(new_n252), .A2(new_n634), .A3(new_n639), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n664), .A2(new_n635), .A3(new_n668), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n590), .A2(new_n591), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n593), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n590), .A2(KEYINPUT73), .A3(new_n591), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n596), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n588), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n679), .A2(G472), .B1(new_n580), .B2(new_n582), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n604), .A2(new_n581), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  INV_X1    g498(.A(new_n584), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n560), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n591), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n567), .A2(new_n568), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n598), .B1(new_n688), .B2(new_n271), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n580), .B2(new_n582), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n690), .A2(new_n691), .A3(new_n681), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n690), .B2(new_n681), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n497), .A2(new_n498), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT38), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n252), .A2(new_n268), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n635), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n654), .A3(new_n624), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n671), .B(KEYINPUT39), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n668), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n700), .B1(KEYINPUT40), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n694), .B(new_n703), .C1(KEYINPUT40), .C2(new_n702), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n618), .A2(new_n615), .A3(new_n613), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n697), .A2(new_n706), .A3(new_n707), .A4(new_n671), .ZN(new_n708));
  INV_X1    g522(.A(G475), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n253), .B1(new_n248), .B2(new_n249), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n223), .A2(new_n249), .A3(new_n233), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n238), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n709), .B1(new_n712), .B2(new_n271), .ZN(new_n713));
  AOI211_X1 g527(.A(KEYINPUT20), .B(new_n637), .C1(new_n238), .C2(new_n259), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n636), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n707), .B(new_n671), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n664), .A2(new_n668), .A3(new_n708), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n682), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  AOI21_X1  g535(.A(new_n545), .B1(new_n680), .B2(new_n681), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n402), .A2(new_n429), .B1(new_n436), .B2(new_n405), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n667), .A3(new_n338), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n625), .A2(new_n725), .A3(new_n619), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n641), .A3(new_n725), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  NOR3_X1   g546(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n725), .A2(KEYINPUT103), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n667), .A3(new_n338), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n735), .B1(new_n736), .B2(new_n663), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n660), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n334), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n738), .B(new_n739), .C1(new_n599), .C2(new_n601), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NOR2_X1   g555(.A1(new_n585), .A2(new_n564), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n571), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n569), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n600), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(new_n546), .C1(new_n598), .C2(new_n606), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n697), .A2(new_n748), .A3(new_n635), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n625), .A3(new_n725), .A4(new_n749), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n734), .A2(new_n737), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n717), .A2(new_n708), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n654), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n745), .B1(new_n598), .B2(new_n606), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n630), .A2(G472), .B1(new_n600), .B2(new_n744), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n738), .A3(KEYINPUT105), .A4(new_n755), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NAND2_X1  g576(.A1(new_n717), .A2(new_n708), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n668), .A2(new_n448), .A3(new_n695), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n722), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT42), .B1(new_n722), .B2(new_n765), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n765), .A2(KEYINPUT42), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n681), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n601), .A2(KEYINPUT107), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n680), .A3(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n779), .A2(KEYINPUT108), .A3(new_n546), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT108), .B1(new_n779), .B2(new_n546), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n197), .ZN(G33));
  NAND2_X1  g598(.A1(new_n672), .A2(new_n635), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n764), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n546), .C1(new_n599), .C2(new_n601), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  NAND2_X1  g602(.A1(new_n695), .A2(new_n448), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n631), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n707), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n697), .A2(KEYINPUT43), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n794), .A2(KEYINPUT43), .B1(new_n707), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n796), .A3(new_n654), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n801), .A3(new_n798), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n801), .B1(new_n797), .B2(new_n798), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n800), .B(KEYINPUT112), .C1(new_n803), .C2(new_n804), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n440), .B1(new_n441), .B2(new_n439), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n443), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n813), .B(new_n814), .C1(new_n810), .C2(new_n809), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n445), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT46), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT46), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n667), .A3(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n819), .A2(new_n338), .A3(new_n701), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n807), .A2(new_n808), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT113), .B(G137), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(G39));
  NOR4_X1   g637(.A1(new_n682), .A2(new_n546), .A3(new_n763), .A4(new_n789), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n819), .A2(KEYINPUT47), .A3(new_n338), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n819), .B2(new_n338), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NOR3_X1   g642(.A1(new_n545), .A2(new_n624), .A3(new_n337), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n724), .A2(new_n667), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OR4_X1    g647(.A1(new_n694), .A2(new_n696), .A3(new_n794), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n825), .A2(new_n826), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n724), .A2(new_n667), .A3(new_n337), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n796), .A2(new_n270), .ZN(new_n838));
  INV_X1    g652(.A(new_n746), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n837), .A2(new_n790), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n694), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n789), .A2(new_n736), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n546), .A3(new_n270), .A4(new_n843), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n844), .A2(new_n697), .A3(new_n707), .ZN(new_n845));
  NAND2_X1  g659(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n846));
  NOR2_X1   g660(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n696), .A2(new_n448), .A3(new_n736), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n838), .A2(new_n843), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n654), .A3(new_n759), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n840), .A2(new_n848), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n849), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n841), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n841), .B2(new_n854), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n844), .A2(new_n620), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n269), .B(new_n858), .C1(new_n754), .C2(new_n840), .ZN(new_n859));
  INV_X1    g673(.A(new_n780), .ZN(new_n860));
  INV_X1    g674(.A(new_n781), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n850), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT48), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n747), .A2(new_n733), .A3(new_n749), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n660), .A2(new_n668), .A3(new_n671), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n692), .B2(new_n693), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n673), .A2(new_n718), .B1(new_n680), .B2(new_n681), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(KEYINPUT114), .A2(new_n761), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n758), .B2(new_n760), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT114), .B1(new_n874), .B2(new_n870), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n866), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n761), .A2(new_n870), .A3(new_n872), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n874), .A2(KEYINPUT114), .A3(new_n870), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n640), .A2(new_n625), .A3(new_n725), .ZN(new_n882));
  AOI221_X4 g696(.A(new_n545), .B1(new_n882), .B2(new_n726), .C1(new_n680), .C2(new_n681), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n713), .A2(new_n715), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n707), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n884), .B2(new_n333), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n500), .A2(new_n502), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n275), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n888), .A2(new_n607), .B1(new_n746), .B2(new_n750), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n740), .A2(new_n602), .A3(new_n655), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n759), .A2(new_n765), .A3(new_n654), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n672), .A2(new_n333), .A3(new_n654), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n764), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n599), .B2(new_n601), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n787), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n890), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n773), .B2(new_n782), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n876), .A2(new_n881), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n877), .A2(KEYINPUT52), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n876), .A2(new_n898), .A3(KEYINPUT53), .A4(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n899), .A2(new_n900), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n876), .A2(new_n898), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n902), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n906), .B(KEYINPUT115), .C1(new_n905), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n901), .A2(new_n903), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n912), .A2(KEYINPUT115), .A3(KEYINPUT54), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n865), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n834), .B1(new_n914), .B2(new_n915), .ZN(G75));
  AOI21_X1  g730(.A(new_n271), .B1(new_n901), .B2(new_n903), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n472), .A2(new_n481), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n479), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n189), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(new_n444), .B(KEYINPUT57), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n904), .A2(new_n905), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n666), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n904), .A2(new_n271), .A3(new_n815), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(G54));
  INV_X1    g747(.A(new_n925), .ZN(new_n934));
  AND2_X1   g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n917), .A2(new_n260), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n260), .B1(new_n917), .B2(new_n935), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n934), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n912), .A2(G902), .A3(new_n935), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n940), .A2(KEYINPUT117), .A3(new_n260), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT118), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT117), .B1(new_n940), .B2(new_n260), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n925), .B1(new_n940), .B2(new_n260), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT118), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n937), .A2(new_n938), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n947), .ZN(G60));
  XOR2_X1   g762(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n949));
  NOR2_X1   g763(.A1(new_n331), .A2(new_n271), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n609), .A2(new_n611), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n928), .B2(new_n929), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n934), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n911), .A2(new_n913), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n609), .A2(new_n611), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(G63));
  INV_X1    g771(.A(KEYINPUT122), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n934), .B1(new_n958), .B2(KEYINPUT61), .ZN(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n277), .A2(new_n271), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n912), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n963), .B2(new_n649), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n912), .A2(new_n962), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n540), .B(KEYINPUT121), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n964), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n964), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n273), .B2(new_n477), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n890), .A2(new_n891), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n920), .B1(G898), .B2(new_n189), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  AND2_X1   g791(.A1(new_n554), .A2(new_n558), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n254), .A2(new_n255), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n702), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n722), .A2(new_n982), .A3(new_n790), .A4(new_n886), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n827), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n704), .A2(new_n874), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n984), .A2(new_n821), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n981), .B1(new_n988), .B2(new_n189), .ZN(new_n989));
  INV_X1    g803(.A(new_n867), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n820), .A2(new_n862), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n827), .A2(new_n991), .A3(new_n787), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(new_n783), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n821), .A2(new_n994), .A3(new_n874), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n821), .B2(new_n874), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n189), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n980), .B1(G900), .B2(G953), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n989), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT124), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n997), .B2(new_n998), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1002), .ZN(new_n1004));
  AOI221_X4 g818(.A(new_n989), .B1(new_n1000), .B2(new_n1004), .C1(new_n997), .C2(new_n998), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(G72));
  OAI211_X1 g820(.A(new_n974), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1007));
  XNOR2_X1  g821(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  AOI211_X1 g824(.A(new_n590), .B(new_n564), .C1(new_n1007), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n974), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1010), .B1(new_n988), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1013), .A2(new_n590), .A3(new_n564), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n595), .A2(new_n567), .A3(new_n568), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1010), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n910), .A2(new_n1016), .ZN(new_n1017));
  NOR4_X1   g831(.A1(new_n1011), .A2(new_n1014), .A3(new_n925), .A4(new_n1017), .ZN(G57));
endmodule


