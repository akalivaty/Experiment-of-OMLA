//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G125), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT16), .A3(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT72), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(KEYINPUT72), .A2(G125), .A3(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n194), .B2(KEYINPUT16), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G237), .ZN(new_n198));
  INV_X1    g012(.A(G953), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G214), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(G237), .A2(G953), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n204), .B(G214), .C1(new_n201), .C2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n197), .B(new_n211), .C1(new_n208), .C2(new_n207), .ZN(new_n212));
  XNOR2_X1  g026(.A(G113), .B(G122), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G125), .B(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n196), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n196), .B2(new_n194), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(new_n209), .ZN(new_n220));
  OAI221_X1 g034(.A(new_n218), .B1(new_n206), .B2(new_n220), .C1(new_n207), .C2(new_n219), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n212), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT93), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT93), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n212), .A2(new_n224), .A3(new_n215), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n212), .A2(new_n221), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n215), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n187), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT20), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n203), .A2(new_n205), .A3(new_n209), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n209), .B1(new_n203), .B2(new_n205), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n207), .A2(KEYINPUT88), .A3(new_n210), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n195), .A2(G146), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n192), .A2(KEYINPUT19), .A3(new_n193), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT89), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT89), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n192), .A2(new_n244), .A3(KEYINPUT19), .A4(new_n193), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n191), .A2(G125), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n188), .A2(G140), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT19), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT90), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n216), .A2(new_n252), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT91), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n246), .A2(new_n254), .A3(new_n255), .A4(new_n196), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n246), .A2(new_n254), .A3(new_n196), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT91), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n239), .A2(new_n241), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n233), .B(new_n215), .C1(new_n259), .C2(new_n221), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n241), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n237), .A2(new_n238), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n221), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n215), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT92), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(G475), .B1(new_n266), .B2(new_n226), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n232), .B1(new_n267), .B2(new_n229), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n233), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n263), .A2(KEYINPUT92), .A3(new_n264), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n226), .A3(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(new_n232), .A3(new_n187), .A4(new_n229), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n231), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n187), .A3(new_n229), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT20), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n273), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT94), .A3(new_n231), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n214), .A2(G107), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n214), .A2(G107), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n288));
  INV_X1    g102(.A(G107), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(G104), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n290), .A3(new_n283), .ZN(new_n291));
  INV_X1    g105(.A(G101), .ZN(new_n292));
  MUX2_X1   g106(.A(new_n286), .B(new_n291), .S(new_n292), .Z(new_n293));
  NAND2_X1  g107(.A1(new_n196), .A2(G143), .ZN(new_n294));
  INV_X1    g108(.A(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G146), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT66), .B(G128), .Z(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(G143), .B2(new_n196), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT64), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n196), .B2(G143), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(KEYINPUT64), .A3(G146), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n299), .A3(G128), .A4(new_n294), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n293), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(KEYINPUT79), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n294), .ZN(new_n310));
  INV_X1    g124(.A(G128), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n300), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n303), .A2(new_n304), .B1(G143), .B2(new_n196), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n299), .A4(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n293), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT80), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n319), .A3(new_n293), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n308), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(G137), .ZN(new_n325));
  INV_X1    g139(.A(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT11), .A3(G134), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G131), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n324), .A2(new_n327), .A3(new_n209), .A4(new_n325), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n321), .A2(KEYINPUT12), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n316), .A2(new_n319), .A3(new_n293), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n319), .B1(new_n316), .B2(new_n293), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n335), .A2(new_n336), .B1(new_n307), .B2(new_n293), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n337), .B2(new_n331), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n335), .B2(new_n336), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n291), .A2(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n291), .A2(KEYINPUT78), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G101), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  INV_X1    g159(.A(new_n291), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(new_n292), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n295), .A2(KEYINPUT64), .A3(G146), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT64), .B1(new_n295), .B2(G146), .ZN(new_n350));
  OAI211_X1 g164(.A(G128), .B(new_n294), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n297), .A2(new_n311), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT0), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n311), .B1(new_n294), .B2(new_n296), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT0), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(G101), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n348), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n293), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n341), .A2(new_n332), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n199), .A2(G227), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n339), .A2(KEYINPUT82), .A3(new_n361), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n318), .B2(new_n320), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n360), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n331), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n361), .A3(KEYINPUT81), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n331), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  INV_X1    g185(.A(new_n364), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT12), .B1(new_n321), .B2(new_n332), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n337), .A2(new_n334), .A3(new_n331), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n374), .A2(new_n361), .A3(new_n375), .A4(new_n364), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n365), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G469), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n229), .ZN(new_n381));
  NAND2_X1  g195(.A1(G469), .A2(G902), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n372), .B1(new_n369), .B2(new_n371), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n374), .A2(new_n361), .A3(new_n375), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n372), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(G469), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT9), .B(G234), .Z(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n229), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(G221), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n391), .B(KEYINPUT77), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G116), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(G122), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n396));
  INV_X1    g210(.A(G122), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(G116), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(KEYINPUT95), .A3(G122), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n289), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n295), .A2(G128), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT66), .B(G128), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n295), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n404), .A2(G134), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n402), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT13), .ZN(new_n407));
  OAI21_X1  g221(.A(G134), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n401), .B(new_n405), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(G134), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT96), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n415));
  OAI21_X1  g229(.A(G107), .B1(new_n395), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n400), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n400), .A2(new_n416), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n389), .A2(G217), .A3(new_n199), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G902), .ZN(new_n425));
  INV_X1    g239(.A(G478), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n426), .A2(KEYINPUT15), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n425), .B(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n282), .A2(new_n393), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT2), .B(G113), .Z(new_n432));
  NOR2_X1   g246(.A1(new_n394), .A2(G119), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT67), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n394), .B2(G119), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n432), .B(new_n434), .C1(new_n433), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(G113), .A3(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT85), .Z(new_n444));
  OAI211_X1 g258(.A(new_n434), .B(KEYINPUT5), .C1(new_n433), .C2(new_n436), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n437), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n293), .ZN(new_n448));
  XOR2_X1   g262(.A(G110), .B(G122), .Z(new_n449));
  XOR2_X1   g263(.A(new_n449), .B(KEYINPUT8), .Z(new_n450));
  OR3_X1    g264(.A1(new_n446), .A2(new_n443), .A3(KEYINPUT84), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT84), .B1(new_n446), .B2(new_n443), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n437), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n448), .B(new_n450), .C1(new_n453), .C2(new_n293), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n199), .A2(G224), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n456));
  AOI21_X1  g270(.A(G128), .B1(new_n294), .B2(new_n296), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n313), .B2(G128), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n355), .B1(new_n458), .B2(KEYINPUT0), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n301), .A2(new_n306), .A3(new_n188), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT86), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(KEYINPUT86), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n456), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n451), .A2(new_n437), .A3(new_n293), .A4(new_n452), .ZN(new_n466));
  INV_X1    g280(.A(new_n449), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n434), .B1(new_n433), .B2(new_n436), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n432), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n348), .A3(new_n358), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n460), .A2(new_n461), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n473), .A2(new_n456), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n454), .A2(new_n465), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n466), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n449), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n473), .B(new_n455), .Z(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n480), .A3(new_n449), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n482), .A3(new_n229), .ZN(new_n483));
  OAI21_X1  g297(.A(G210), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n475), .A2(new_n482), .A3(new_n229), .A4(new_n484), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n431), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(KEYINPUT97), .A2(G952), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT97), .A2(G952), .ZN(new_n491));
  AOI21_X1  g305(.A(G953), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G234), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n493), .B2(new_n198), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT21), .B(G898), .Z(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n229), .B(new_n199), .C1(G234), .C2(G237), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n429), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G217), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(G234), .B2(new_n229), .ZN(new_n503));
  INV_X1    g317(.A(new_n197), .ZN(new_n504));
  INV_X1    g318(.A(G119), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n403), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT71), .B(KEYINPUT23), .Z(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n505), .B2(G128), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n507), .B(new_n509), .C1(G119), .C2(new_n311), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G110), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n506), .B1(new_n505), .B2(G128), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT24), .B(G110), .Z(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n504), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n504), .A2(new_n511), .A3(new_n517), .A4(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n510), .A2(G110), .B1(new_n512), .B2(new_n513), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  OAI221_X1 g336(.A(new_n522), .B1(new_n512), .B2(new_n513), .C1(new_n510), .C2(G110), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n521), .A2(new_n241), .A3(new_n523), .A4(new_n217), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n199), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(new_n524), .A3(new_n530), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT25), .B1(new_n534), .B2(new_n229), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n519), .A2(new_n524), .A3(new_n530), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n519), .B2(new_n524), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT25), .B(new_n229), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n503), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n503), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(G472), .A2(G902), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n326), .A2(G134), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n323), .A2(G137), .ZN(new_n548));
  OAI21_X1  g362(.A(G131), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n330), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n307), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT30), .B(new_n551), .C1(new_n459), .C2(new_n332), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT65), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n330), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n330), .B2(new_n549), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n556), .A2(new_n307), .B1(new_n357), .B2(new_n331), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n470), .B(new_n552), .C1(new_n557), .C2(KEYINPUT30), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n357), .A2(new_n331), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n469), .A3(new_n551), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n198), .A2(new_n199), .A3(G210), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT27), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT26), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n292), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n563), .B(KEYINPUT26), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G101), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n558), .A2(new_n560), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT68), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n558), .A2(KEYINPUT68), .A3(new_n560), .A4(new_n569), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n546), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n557), .A2(new_n469), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n568), .ZN(new_n579));
  INV_X1    g393(.A(new_n566), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT69), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT69), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n566), .B2(new_n568), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n578), .A2(new_n584), .B1(new_n570), .B2(KEYINPUT31), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n545), .B1(new_n574), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(KEYINPUT70), .B(new_n545), .C1(new_n574), .C2(new_n585), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT32), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n569), .B1(new_n558), .B2(new_n560), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT29), .B(new_n591), .C1(new_n578), .C2(new_n584), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n559), .A2(new_n551), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n470), .ZN(new_n594));
  INV_X1    g408(.A(new_n577), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n569), .A2(KEYINPUT29), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n229), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G472), .B1(new_n592), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT32), .B(new_n545), .C1(new_n574), .C2(new_n585), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n590), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n544), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n501), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  INV_X1    g420(.A(new_n393), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n588), .A2(new_n589), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n229), .B1(new_n574), .B2(new_n585), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n607), .A2(new_n608), .A3(new_n543), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n543), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT98), .B1(new_n615), .B2(new_n393), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n422), .B2(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n424), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n424), .ZN(new_n621));
  OAI211_X1 g435(.A(G478), .B(new_n229), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n426), .B1(new_n424), .B2(G902), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n277), .B2(new_n281), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n500), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(KEYINPUT100), .A3(new_n500), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n617), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT101), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT34), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n214), .ZN(G6));
  NAND3_X1  g447(.A1(new_n279), .A2(KEYINPUT102), .A3(new_n273), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT102), .B1(new_n279), .B2(new_n273), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n428), .B(new_n231), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n637), .A2(new_n499), .A3(new_n489), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NOR2_X1   g455(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n525), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n541), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n612), .B1(new_n540), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n501), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT37), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G110), .ZN(G12));
  INV_X1    g462(.A(new_n636), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n634), .ZN(new_n650));
  INV_X1    g464(.A(new_n498), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(G900), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n494), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n650), .A2(new_n428), .A3(new_n231), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n540), .A2(new_n644), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n655), .B(new_n488), .C1(new_n590), .C2(new_n602), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n654), .A2(new_n656), .A3(new_n393), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n656), .A2(new_n393), .ZN(new_n659));
  INV_X1    g473(.A(new_n653), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n637), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT104), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n311), .ZN(G30));
  INV_X1    g478(.A(new_n428), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n277), .B2(new_n281), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n486), .A2(new_n487), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT38), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n430), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n653), .B(KEYINPUT39), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n607), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n601), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  INV_X1    g489(.A(new_n584), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n594), .A2(new_n560), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n572), .A2(new_n573), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n676), .A2(KEYINPUT105), .A3(new_n677), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n675), .B1(new_n683), .B2(new_n229), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n590), .A2(new_n674), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n655), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n673), .B(new_n686), .C1(new_n672), .C2(new_n671), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NAND2_X1  g502(.A1(new_n622), .A2(new_n623), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT94), .B1(new_n280), .B2(new_n231), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n276), .B(new_n230), .C1(new_n279), .C2(new_n273), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n689), .B(new_n653), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n659), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  AND3_X1   g509(.A1(new_n379), .A2(new_n380), .A3(new_n229), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n380), .B1(new_n379), .B2(new_n229), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n696), .A2(new_n697), .A3(new_n391), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n699), .A2(new_n603), .A3(new_n544), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n628), .A2(new_n629), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n638), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND2_X1  g519(.A1(new_n379), .A2(new_n229), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  INV_X1    g521(.A(new_n391), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n488), .A3(new_n381), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n282), .A2(new_n603), .A3(new_n499), .A4(new_n428), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n655), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NAND4_X1  g528(.A1(new_n282), .A2(KEYINPUT108), .A3(new_n488), .A4(new_n428), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n488), .B(new_n428), .C1(new_n690), .C2(new_n691), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n597), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n597), .A2(new_n720), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n676), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n574), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n723), .B(new_n724), .C1(KEYINPUT31), .C2(new_n570), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n725), .A2(new_n545), .B1(G472), .B2(new_n610), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n543), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n699), .A2(new_n727), .A3(new_n499), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  AND2_X1   g544(.A1(new_n726), .A2(new_n655), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT106), .B1(new_n698), .B2(new_n488), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n709), .A2(new_n710), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n731), .B(new_n693), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  XNOR2_X1  g549(.A(new_n382), .B(KEYINPUT109), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n381), .A2(new_n387), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT110), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n486), .A2(new_n430), .A3(new_n487), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n391), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n693), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT32), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n586), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n602), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n544), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT42), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n738), .A3(new_n604), .A4(new_n740), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n209), .ZN(G33));
  NAND4_X1  g565(.A1(new_n738), .A2(new_n661), .A3(new_n604), .A4(new_n740), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NAND3_X1  g567(.A1(new_n384), .A2(KEYINPUT45), .A3(new_n386), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  INV_X1    g569(.A(new_n386), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n383), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n757), .A3(G469), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT46), .A3(new_n736), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n381), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT111), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n736), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(new_n765), .A3(new_n381), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n761), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n708), .A3(new_n670), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT112), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n739), .B(KEYINPUT114), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT113), .B1(new_n282), .B2(new_n624), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT113), .B(KEYINPUT43), .C1(new_n282), .C2(new_n624), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n612), .A3(new_n655), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n770), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n769), .B(new_n777), .C1(new_n776), .C2(new_n775), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  NAND2_X1  g593(.A1(new_n767), .A2(new_n708), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n692), .A2(new_n543), .A3(new_n739), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n767), .A2(new_n783), .A3(new_n708), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n603), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n685), .A2(new_n391), .A3(new_n655), .A4(new_n660), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT108), .B1(new_n666), .B2(new_n488), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n716), .A2(new_n717), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n788), .B(new_n738), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n737), .B(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n718), .B2(new_n715), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT115), .A3(new_n788), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n734), .B(new_n694), .C1(new_n658), .C2(new_n662), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n787), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n799), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT52), .A3(new_n793), .A4(new_n797), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n734), .B1(new_n658), .B2(new_n662), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n701), .A2(new_n713), .A3(new_n704), .A4(new_n729), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n282), .A2(new_n689), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n665), .B2(new_n282), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n614), .A3(new_n616), .A4(new_n500), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n429), .B(new_n500), .C1(new_n604), .C2(new_n645), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n739), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n655), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n603), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n660), .B(new_n428), .C1(new_n649), .C2(new_n634), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n607), .A4(new_n231), .ZN(new_n818));
  INV_X1    g632(.A(new_n731), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n752), .B(new_n818), .C1(new_n741), .C2(new_n819), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n808), .A2(new_n750), .A3(new_n813), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n803), .A2(new_n807), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT53), .B1(new_n803), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n791), .A2(new_n792), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n796), .B2(new_n788), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(new_n827), .B2(new_n801), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n798), .A2(new_n787), .A3(new_n799), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n821), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n806), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n806), .B1(new_n804), .B2(KEYINPUT52), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n803), .A2(new_n821), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n696), .A2(new_n697), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(new_n740), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n543), .A2(new_n839), .A3(new_n495), .A4(new_n685), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n625), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n773), .A2(new_n495), .A3(new_n774), .A4(new_n839), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n746), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT48), .Z(new_n844));
  INV_X1    g658(.A(new_n727), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n773), .A2(new_n495), .A3(new_n845), .A4(new_n774), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n711), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n492), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n282), .A2(new_n689), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n840), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n842), .B2(new_n819), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n392), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n781), .A2(new_n784), .B1(new_n855), .B2(new_n838), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n846), .A2(new_n770), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n854), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n850), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n781), .A2(new_n784), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n838), .A2(new_n855), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n853), .B1(new_n864), .B2(new_n857), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n668), .A2(new_n430), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n847), .A2(new_n698), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT50), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n847), .A2(KEYINPUT50), .A3(new_n698), .A4(new_n866), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n865), .A2(new_n871), .A3(new_n860), .A4(new_n850), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n849), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n836), .A2(new_n837), .A3(new_n841), .A4(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(G952), .A2(G953), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n824), .A3(new_n835), .A4(new_n841), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n668), .A2(new_n855), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n881), .A2(new_n430), .A3(new_n685), .ZN(new_n882));
  INV_X1    g696(.A(new_n838), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n624), .B(new_n282), .C1(KEYINPUT49), .C2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(KEYINPUT49), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n884), .A3(new_n543), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n886), .ZN(G75));
  AND3_X1   g701(.A1(new_n803), .A2(new_n821), .A3(new_n833), .ZN(new_n888));
  OAI211_X1 g702(.A(G210), .B(G902), .C1(new_n888), .C2(new_n823), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT119), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n892), .A3(new_n890), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n478), .A2(new_n481), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n479), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  AOI22_X1  g710(.A1(KEYINPUT118), .A2(new_n891), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n891), .A2(KEYINPUT118), .A3(new_n896), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n199), .A2(G952), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G51));
  OAI21_X1  g714(.A(KEYINPUT54), .B1(new_n888), .B2(new_n823), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n835), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n736), .B(KEYINPUT57), .Z(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n379), .B(KEYINPUT120), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n229), .B1(new_n831), .B2(new_n834), .ZN(new_n907));
  INV_X1    g721(.A(new_n758), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n906), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  INV_X1    g725(.A(new_n272), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n899), .ZN(G60));
  OR2_X1    g729(.A1(new_n620), .A2(new_n621), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n824), .A2(new_n835), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n916), .A2(new_n920), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n899), .B(new_n921), .C1(new_n902), .C2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT123), .Z(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT60), .Z(new_n926));
  OAI211_X1 g740(.A(new_n643), .B(new_n926), .C1(new_n888), .C2(new_n823), .ZN(new_n927));
  INV_X1    g741(.A(new_n899), .ZN(new_n928));
  INV_X1    g742(.A(new_n926), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n831), .B2(new_n834), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n927), .B(new_n928), .C1(new_n930), .C2(new_n534), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT122), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT61), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT124), .B1(new_n931), .B2(KEYINPUT122), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n931), .B2(KEYINPUT124), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n934), .B1(new_n935), .B2(new_n937), .ZN(G66));
  AOI21_X1  g752(.A(new_n199), .B1(new_n496), .B2(G224), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n808), .A2(new_n813), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n199), .ZN(new_n941));
  MUX2_X1   g755(.A(new_n939), .B(new_n941), .S(KEYINPUT125), .Z(new_n942));
  INV_X1    g756(.A(G898), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n894), .B1(new_n943), .B2(G953), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G69));
  OAI21_X1  g759(.A(new_n552), .B1(new_n557), .B2(KEYINPUT30), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n246), .A2(new_n254), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT126), .Z(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(G900), .B1(new_n950), .B2(G227), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n199), .B(new_n951), .C1(G227), .C2(new_n950), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n778), .A2(new_n785), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n769), .A2(new_n719), .A3(new_n745), .ZN(new_n954));
  INV_X1    g768(.A(new_n752), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n750), .A2(new_n799), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(new_n949), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n810), .A2(new_n671), .A3(new_n604), .A4(new_n814), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n801), .A2(new_n687), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT62), .Z(new_n961));
  NAND3_X1  g775(.A1(new_n953), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(G953), .B1(new_n962), .B2(new_n949), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(new_n958), .B2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n957), .B2(new_n940), .ZN(new_n967));
  INV_X1    g781(.A(new_n569), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n560), .A3(new_n558), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n966), .B1(new_n962), .B2(new_n940), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n558), .A2(new_n560), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n971), .A3(new_n569), .ZN(new_n972));
  INV_X1    g786(.A(new_n966), .ZN(new_n973));
  INV_X1    g787(.A(new_n591), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n681), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n822), .B2(new_n823), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n928), .A2(new_n969), .A3(new_n972), .A4(new_n977), .ZN(G57));
endmodule


