

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709;

  XNOR2_X2 U363 ( .A(n339), .B(n568), .ZN(n683) );
  NAND2_X1 U364 ( .A1(n567), .A2(n346), .ZN(n339) );
  XNOR2_X1 U365 ( .A(n349), .B(G119), .ZN(n436) );
  NOR2_X1 U366 ( .A1(n498), .A2(n497), .ZN(n351) );
  INV_X1 U367 ( .A(G953), .ZN(n700) );
  NOR2_X1 U368 ( .A1(n361), .A2(n557), .ZN(n564) );
  XNOR2_X1 U369 ( .A(n552), .B(KEYINPUT35), .ZN(n361) );
  XNOR2_X1 U370 ( .A(n532), .B(n531), .ZN(n352) );
  NOR2_X1 U371 ( .A1(n487), .A2(n469), .ZN(n471) );
  XNOR2_X1 U372 ( .A(n351), .B(n348), .ZN(n527) );
  XNOR2_X1 U373 ( .A(n363), .B(n342), .ZN(n675) );
  NOR2_X1 U374 ( .A1(G902), .A2(n665), .ZN(n410) );
  XNOR2_X1 U375 ( .A(KEYINPUT66), .B(KEYINPUT83), .ZN(n396) );
  XNOR2_X2 U376 ( .A(n350), .B(n528), .ZN(n539) );
  XNOR2_X1 U377 ( .A(n401), .B(n400), .ZN(n457) );
  NOR2_X1 U378 ( .A1(n709), .A2(n705), .ZN(n485) );
  XNOR2_X1 U379 ( .A(n402), .B(G134), .ZN(n369) );
  XOR2_X1 U380 ( .A(G137), .B(G131), .Z(n402) );
  XNOR2_X1 U381 ( .A(n617), .B(KEYINPUT86), .ZN(n366) );
  AND2_X1 U382 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U383 ( .A(n376), .B(n375), .ZN(n692) );
  XNOR2_X1 U384 ( .A(G125), .B(G140), .ZN(n375) );
  XOR2_X1 U385 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n376) );
  XNOR2_X1 U386 ( .A(n498), .B(KEYINPUT38), .ZN(n592) );
  XNOR2_X1 U387 ( .A(n478), .B(KEYINPUT41), .ZN(n608) );
  NOR2_X1 U388 ( .A1(n595), .A2(n594), .ZN(n478) );
  XNOR2_X1 U389 ( .A(n362), .B(n425), .ZN(n427) );
  XNOR2_X1 U390 ( .A(n461), .B(n407), .ZN(n408) );
  INV_X1 U391 ( .A(G140), .ZN(n405) );
  AND2_X1 U392 ( .A1(n628), .A2(G953), .ZN(n678) );
  XNOR2_X1 U393 ( .A(n663), .B(KEYINPUT88), .ZN(n367) );
  XNOR2_X1 U394 ( .A(n365), .B(KEYINPUT85), .ZN(n364) );
  NAND2_X1 U395 ( .A1(n366), .A2(n492), .ZN(n365) );
  INV_X1 U396 ( .A(KEYINPUT44), .ZN(n565) );
  XNOR2_X1 U397 ( .A(n474), .B(n473), .ZN(n595) );
  INV_X1 U398 ( .A(KEYINPUT111), .ZN(n473) );
  AND2_X1 U399 ( .A1(n494), .A2(n476), .ZN(n356) );
  AND2_X1 U400 ( .A1(n553), .A2(n357), .ZN(n494) );
  AND2_X1 U401 ( .A1(n358), .A2(n578), .ZN(n357) );
  INV_X1 U402 ( .A(n479), .ZN(n358) );
  XNOR2_X1 U403 ( .A(n475), .B(n360), .ZN(n491) );
  INV_X1 U404 ( .A(n491), .ZN(n359) );
  XNOR2_X1 U405 ( .A(n693), .B(n442), .ZN(n638) );
  XNOR2_X1 U406 ( .A(G107), .B(G116), .ZN(n392) );
  XNOR2_X1 U407 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n470) );
  NAND2_X1 U408 ( .A1(n352), .A2(n543), .ZN(n560) );
  INV_X1 U409 ( .A(KEYINPUT0), .ZN(n528) );
  XNOR2_X1 U410 ( .A(n560), .B(KEYINPUT89), .ZN(n534) );
  INV_X1 U411 ( .A(n535), .ZN(n533) );
  XNOR2_X1 U412 ( .A(n423), .B(n422), .ZN(n363) );
  NOR2_X1 U413 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U414 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n483) );
  NOR2_X1 U415 ( .A1(n608), .A2(n501), .ZN(n484) );
  NAND2_X1 U416 ( .A1(n353), .A2(n579), .ZN(n619) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n353) );
  INV_X1 U418 ( .A(KEYINPUT90), .ZN(n354) );
  NAND2_X1 U419 ( .A1(n534), .A2(n533), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X1 U421 ( .A1(n540), .A2(n546), .ZN(n340) );
  XOR2_X1 U422 ( .A(n440), .B(n439), .Z(n341) );
  XNOR2_X1 U423 ( .A(G146), .B(n692), .ZN(n342) );
  XOR2_X1 U424 ( .A(G128), .B(G143), .Z(n343) );
  XOR2_X1 U425 ( .A(KEYINPUT65), .B(KEYINPUT4), .Z(n344) );
  AND2_X1 U426 ( .A1(n356), .A2(n359), .ZN(n345) );
  AND2_X1 U427 ( .A1(n619), .A2(n542), .ZN(n346) );
  AND2_X1 U428 ( .A1(n493), .A2(n345), .ZN(n347) );
  XOR2_X1 U429 ( .A(n499), .B(KEYINPUT19), .Z(n348) );
  XNOR2_X2 U430 ( .A(G116), .B(KEYINPUT3), .ZN(n349) );
  NAND2_X1 U431 ( .A1(n527), .A2(n526), .ZN(n350) );
  NAND2_X1 U432 ( .A1(n352), .A2(n556), .ZN(n652) );
  NAND2_X1 U433 ( .A1(n359), .A2(n476), .ZN(n644) );
  INV_X1 U434 ( .A(KEYINPUT103), .ZN(n360) );
  XNOR2_X1 U435 ( .A(n361), .B(G122), .ZN(n706) );
  NOR2_X1 U436 ( .A1(n675), .A2(G902), .ZN(n362) );
  NAND2_X1 U437 ( .A1(n367), .A2(n364), .ZN(n507) );
  NAND2_X1 U438 ( .A1(n368), .A2(n535), .ZN(n663) );
  XNOR2_X1 U439 ( .A(n495), .B(KEYINPUT36), .ZN(n368) );
  XNOR2_X2 U440 ( .A(n457), .B(n369), .ZN(n693) );
  BUF_X1 U441 ( .A(n620), .Z(n574) );
  NAND2_X1 U442 ( .A1(n592), .A2(n591), .ZN(n474) );
  INV_X1 U443 ( .A(n592), .ZN(n469) );
  XNOR2_X1 U444 ( .A(n471), .B(n470), .ZN(n511) );
  XNOR2_X1 U445 ( .A(n693), .B(n408), .ZN(n665) );
  XOR2_X1 U446 ( .A(KEYINPUT53), .B(n615), .Z(G75) );
  XOR2_X1 U447 ( .A(KEYINPUT51), .B(n590), .Z(n371) );
  AND2_X1 U448 ( .A1(n506), .A2(n505), .ZN(n372) );
  NOR2_X1 U449 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U450 ( .A1(n507), .A2(n372), .ZN(n508) );
  NOR2_X1 U451 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U452 ( .A(n441), .B(n341), .ZN(n442) );
  XNOR2_X1 U453 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U454 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U455 ( .A(n484), .B(n483), .ZN(n705) );
  XOR2_X1 U456 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n374) );
  XNOR2_X1 U457 ( .A(KEYINPUT13), .B(G475), .ZN(n373) );
  XNOR2_X1 U458 ( .A(n374), .B(n373), .ZN(n388) );
  XOR2_X1 U459 ( .A(KEYINPUT99), .B(G113), .Z(n378) );
  XNOR2_X1 U460 ( .A(G122), .B(G104), .ZN(n377) );
  XNOR2_X1 U461 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U462 ( .A(n342), .B(n379), .Z(n386) );
  XOR2_X1 U463 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n381) );
  NOR2_X1 U464 ( .A1(G953), .A2(G237), .ZN(n437) );
  NAND2_X1 U465 ( .A1(n437), .A2(G214), .ZN(n380) );
  XNOR2_X1 U466 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U467 ( .A(n382), .B(KEYINPUT100), .Z(n384) );
  XNOR2_X1 U468 ( .A(G143), .B(G131), .ZN(n383) );
  XNOR2_X1 U469 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U470 ( .A(n386), .B(n385), .ZN(n670) );
  NOR2_X1 U471 ( .A1(G902), .A2(n670), .ZN(n387) );
  XNOR2_X1 U472 ( .A(n388), .B(n387), .ZN(n486) );
  INV_X1 U473 ( .A(n486), .ZN(n475) );
  NAND2_X1 U474 ( .A1(G234), .A2(n700), .ZN(n389) );
  XOR2_X1 U475 ( .A(KEYINPUT8), .B(n389), .Z(n421) );
  NAND2_X1 U476 ( .A1(G217), .A2(n421), .ZN(n391) );
  XOR2_X1 U477 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n390) );
  XNOR2_X1 U478 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U479 ( .A(G134), .B(G122), .Z(n393) );
  XNOR2_X1 U480 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U481 ( .A(n395), .B(n394), .ZN(n397) );
  XNOR2_X1 U482 ( .A(n343), .B(n396), .ZN(n400) );
  XNOR2_X1 U483 ( .A(n397), .B(n400), .ZN(n632) );
  NOR2_X1 U484 ( .A1(n632), .A2(G902), .ZN(n398) );
  XOR2_X1 U485 ( .A(G478), .B(n398), .Z(n490) );
  INV_X1 U486 ( .A(n490), .ZN(n476) );
  XNOR2_X1 U487 ( .A(KEYINPUT68), .B(G146), .ZN(n399) );
  XOR2_X1 U488 ( .A(n344), .B(n399), .Z(n401) );
  XOR2_X1 U489 ( .A(G101), .B(G104), .Z(n404) );
  XNOR2_X1 U490 ( .A(G107), .B(G110), .ZN(n403) );
  XNOR2_X1 U491 ( .A(n404), .B(n403), .ZN(n679) );
  XNOR2_X1 U492 ( .A(n679), .B(KEYINPUT71), .ZN(n461) );
  NAND2_X1 U493 ( .A1(G227), .A2(n700), .ZN(n406) );
  INV_X1 U494 ( .A(G469), .ZN(n409) );
  XNOR2_X2 U495 ( .A(n410), .B(n409), .ZN(n496) );
  XNOR2_X1 U496 ( .A(KEYINPUT15), .B(G902), .ZN(n621) );
  NAND2_X1 U497 ( .A1(n621), .A2(G234), .ZN(n412) );
  XNOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT98), .ZN(n411) );
  XNOR2_X1 U499 ( .A(n412), .B(n411), .ZN(n424) );
  NAND2_X1 U500 ( .A1(n424), .A2(G221), .ZN(n414) );
  INV_X1 U501 ( .A(KEYINPUT21), .ZN(n413) );
  XNOR2_X1 U502 ( .A(n414), .B(n413), .ZN(n578) );
  INV_X1 U503 ( .A(n578), .ZN(n529) );
  XOR2_X1 U504 ( .A(G137), .B(G119), .Z(n416) );
  XNOR2_X1 U505 ( .A(G128), .B(G110), .ZN(n415) );
  XNOR2_X1 U506 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U507 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n418) );
  XNOR2_X1 U508 ( .A(KEYINPUT96), .B(KEYINPUT24), .ZN(n417) );
  XNOR2_X1 U509 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U510 ( .A(n420), .B(n419), .Z(n423) );
  NAND2_X1 U511 ( .A1(G221), .A2(n421), .ZN(n422) );
  NAND2_X1 U512 ( .A1(G217), .A2(n424), .ZN(n425) );
  XOR2_X1 U513 ( .A(KEYINPUT78), .B(KEYINPUT25), .Z(n426) );
  XNOR2_X1 U514 ( .A(n427), .B(n426), .ZN(n553) );
  NOR2_X1 U515 ( .A1(n529), .A2(n553), .ZN(n583) );
  NAND2_X1 U516 ( .A1(n496), .A2(n583), .ZN(n538) );
  XNOR2_X1 U517 ( .A(KEYINPUT109), .B(n538), .ZN(n449) );
  NAND2_X1 U518 ( .A1(G237), .A2(G234), .ZN(n428) );
  XNOR2_X1 U519 ( .A(KEYINPUT14), .B(n428), .ZN(n431) );
  AND2_X1 U520 ( .A1(G953), .A2(n431), .ZN(n429) );
  NAND2_X1 U521 ( .A1(G902), .A2(n429), .ZN(n523) );
  XNOR2_X1 U522 ( .A(KEYINPUT106), .B(n523), .ZN(n430) );
  NOR2_X1 U523 ( .A1(G900), .A2(n430), .ZN(n433) );
  NAND2_X1 U524 ( .A1(n431), .A2(G952), .ZN(n432) );
  XOR2_X1 U525 ( .A(KEYINPUT95), .B(n432), .Z(n605) );
  NOR2_X1 U526 ( .A1(n605), .A2(G953), .ZN(n522) );
  NOR2_X1 U527 ( .A1(n433), .A2(n522), .ZN(n479) );
  INV_X1 U528 ( .A(KEYINPUT70), .ZN(n434) );
  XNOR2_X1 U529 ( .A(n434), .B(G113), .ZN(n435) );
  XNOR2_X2 U530 ( .A(n436), .B(n435), .ZN(n460) );
  AND2_X1 U531 ( .A1(n437), .A2(G210), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n460), .B(n438), .ZN(n441) );
  XOR2_X1 U533 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n440) );
  XNOR2_X1 U534 ( .A(G101), .B(KEYINPUT5), .ZN(n439) );
  INV_X1 U535 ( .A(G902), .ZN(n445) );
  NAND2_X1 U536 ( .A1(n638), .A2(n445), .ZN(n443) );
  XNOR2_X2 U537 ( .A(n443), .B(G472), .ZN(n577) );
  INV_X1 U538 ( .A(G237), .ZN(n444) );
  NAND2_X1 U539 ( .A1(n445), .A2(n444), .ZN(n465) );
  NAND2_X1 U540 ( .A1(n465), .A2(G214), .ZN(n591) );
  NAND2_X1 U541 ( .A1(n577), .A2(n591), .ZN(n446) );
  XNOR2_X1 U542 ( .A(KEYINPUT30), .B(n446), .ZN(n447) );
  NOR2_X1 U543 ( .A1(n479), .A2(n447), .ZN(n448) );
  NAND2_X1 U544 ( .A1(n449), .A2(n448), .ZN(n487) );
  XOR2_X1 U545 ( .A(KEYINPUT93), .B(G125), .Z(n451) );
  XOR2_X1 U546 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n450) );
  XNOR2_X1 U547 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U548 ( .A(KEYINPUT92), .B(KEYINPUT79), .ZN(n453) );
  NAND2_X1 U549 ( .A1(G224), .A2(n700), .ZN(n452) );
  XNOR2_X1 U550 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U552 ( .A(n457), .B(n456), .ZN(n463) );
  XNOR2_X1 U553 ( .A(KEYINPUT16), .B(G122), .ZN(n458) );
  XNOR2_X1 U554 ( .A(n458), .B(KEYINPUT74), .ZN(n459) );
  XNOR2_X2 U555 ( .A(n460), .B(n459), .ZN(n680) );
  XNOR2_X1 U556 ( .A(n680), .B(n461), .ZN(n462) );
  XNOR2_X1 U557 ( .A(n463), .B(n462), .ZN(n625) );
  INV_X1 U558 ( .A(n621), .ZN(n464) );
  OR2_X2 U559 ( .A1(n625), .A2(n464), .ZN(n468) );
  NAND2_X1 U560 ( .A1(n465), .A2(G210), .ZN(n466) );
  XNOR2_X1 U561 ( .A(n466), .B(KEYINPUT94), .ZN(n467) );
  XNOR2_X2 U562 ( .A(n468), .B(n467), .ZN(n498) );
  NOR2_X1 U563 ( .A1(n644), .A2(n511), .ZN(n472) );
  XNOR2_X1 U564 ( .A(n472), .B(KEYINPUT40), .ZN(n709) );
  NAND2_X1 U565 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U566 ( .A(n477), .B(KEYINPUT104), .ZN(n594) );
  XOR2_X1 U567 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n481) );
  NAND2_X1 U568 ( .A1(n577), .A2(n494), .ZN(n480) );
  XNOR2_X1 U569 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U570 ( .A1(n482), .A2(n496), .ZN(n501) );
  XNOR2_X1 U571 ( .A(n485), .B(KEYINPUT46), .ZN(n509) );
  NAND2_X1 U572 ( .A1(n486), .A2(n490), .ZN(n549) );
  NOR2_X1 U573 ( .A1(n487), .A2(n549), .ZN(n489) );
  INV_X1 U574 ( .A(n498), .ZN(n488) );
  NAND2_X1 U575 ( .A1(n489), .A2(n488), .ZN(n617) );
  NAND2_X1 U576 ( .A1(n491), .A2(n490), .ZN(n647) );
  AND2_X1 U577 ( .A1(n644), .A2(n647), .ZN(n596) );
  NAND2_X1 U578 ( .A1(KEYINPUT47), .A2(n596), .ZN(n492) );
  XNOR2_X1 U579 ( .A(n577), .B(KEYINPUT6), .ZN(n543) );
  INV_X1 U580 ( .A(n543), .ZN(n493) );
  NAND2_X1 U581 ( .A1(n347), .A2(n591), .ZN(n513) );
  NOR2_X1 U582 ( .A1(n513), .A2(n498), .ZN(n495) );
  XNOR2_X2 U583 ( .A(n496), .B(KEYINPUT1), .ZN(n535) );
  INV_X1 U584 ( .A(n591), .ZN(n497) );
  INV_X1 U585 ( .A(KEYINPUT77), .ZN(n499) );
  INV_X1 U586 ( .A(n527), .ZN(n500) );
  NOR2_X1 U587 ( .A1(n501), .A2(n500), .ZN(n655) );
  NAND2_X1 U588 ( .A1(n644), .A2(n647), .ZN(n502) );
  NAND2_X1 U589 ( .A1(n655), .A2(n502), .ZN(n504) );
  INV_X1 U590 ( .A(KEYINPUT47), .ZN(n503) );
  NAND2_X1 U591 ( .A1(n504), .A2(n503), .ZN(n506) );
  NAND2_X1 U592 ( .A1(n655), .A2(KEYINPUT47), .ZN(n505) );
  XNOR2_X1 U593 ( .A(n510), .B(KEYINPUT48), .ZN(n521) );
  OR2_X1 U594 ( .A1(n511), .A2(n647), .ZN(n512) );
  XNOR2_X1 U595 ( .A(n512), .B(KEYINPUT113), .ZN(n704) );
  NOR2_X1 U596 ( .A1(n535), .A2(n513), .ZN(n515) );
  XNOR2_X1 U597 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U598 ( .A(n515), .B(n514), .ZN(n516) );
  AND2_X1 U599 ( .A1(n516), .A2(n498), .ZN(n518) );
  INV_X1 U600 ( .A(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U601 ( .A(n518), .B(n517), .ZN(n707) );
  INV_X1 U602 ( .A(n707), .ZN(n519) );
  NOR2_X1 U603 ( .A1(n704), .A2(n519), .ZN(n520) );
  NAND2_X1 U604 ( .A1(n521), .A2(n520), .ZN(n698) );
  INV_X1 U605 ( .A(n522), .ZN(n525) );
  OR2_X1 U606 ( .A1(n523), .A2(G898), .ZN(n524) );
  NAND2_X1 U607 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U608 ( .A1(n594), .A2(n529), .ZN(n530) );
  NAND2_X1 U609 ( .A1(n539), .A2(n530), .ZN(n532) );
  XNOR2_X1 U610 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n531) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT105), .ZN(n579) );
  NAND2_X1 U612 ( .A1(n583), .A2(n535), .ZN(n544) );
  INV_X1 U613 ( .A(n544), .ZN(n536) );
  AND2_X1 U614 ( .A1(n577), .A2(n536), .ZN(n589) );
  NAND2_X1 U615 ( .A1(n539), .A2(n589), .ZN(n537) );
  XNOR2_X1 U616 ( .A(n537), .B(KEYINPUT31), .ZN(n660) );
  OR2_X1 U617 ( .A1(n538), .A2(n577), .ZN(n540) );
  INV_X1 U618 ( .A(n539), .ZN(n546) );
  NOR2_X1 U619 ( .A1(n660), .A2(n340), .ZN(n541) );
  OR2_X1 U620 ( .A1(n541), .A2(n596), .ZN(n542) );
  XNOR2_X1 U621 ( .A(n545), .B(KEYINPUT33), .ZN(n599) );
  NOR2_X1 U622 ( .A1(n599), .A2(n546), .ZN(n548) );
  XOR2_X1 U623 ( .A(KEYINPUT34), .B(KEYINPUT81), .Z(n547) );
  XNOR2_X1 U624 ( .A(n548), .B(n547), .ZN(n551) );
  XOR2_X1 U625 ( .A(n549), .B(KEYINPUT80), .Z(n550) );
  NAND2_X1 U626 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U627 ( .A(n553), .ZN(n554) );
  OR2_X1 U628 ( .A1(n577), .A2(n554), .ZN(n555) );
  NOR2_X1 U629 ( .A1(n535), .A2(n555), .ZN(n556) );
  INV_X1 U630 ( .A(n652), .ZN(n557) );
  INV_X1 U631 ( .A(n579), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n535), .A2(n558), .ZN(n559) );
  NOR2_X1 U633 ( .A1(n560), .A2(n559), .ZN(n563) );
  XNOR2_X1 U634 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n561) );
  XNOR2_X1 U635 ( .A(n561), .B(KEYINPUT67), .ZN(n562) );
  XNOR2_X1 U636 ( .A(n563), .B(n562), .ZN(n618) );
  NAND2_X1 U637 ( .A1(n564), .A2(n618), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U639 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n568) );
  NOR2_X2 U640 ( .A1(n698), .A2(n683), .ZN(n620) );
  INV_X1 U641 ( .A(n574), .ZN(n571) );
  XOR2_X1 U642 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n570) );
  NAND2_X1 U643 ( .A1(n571), .A2(n570), .ZN(n576) );
  INV_X1 U644 ( .A(KEYINPUT2), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n572), .A2(KEYINPUT84), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n613) );
  INV_X1 U648 ( .A(n577), .ZN(n582) );
  NOR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT49), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n586) );
  NOR2_X1 U652 ( .A1(n583), .A2(n535), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT50), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT119), .B(n587), .Z(n588) );
  NOR2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n608), .A2(n371), .ZN(n602) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n598) );
  NOR2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n600) );
  NOR2_X1 U661 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U662 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U663 ( .A(KEYINPUT52), .B(n603), .ZN(n604) );
  XOR2_X1 U664 ( .A(KEYINPUT120), .B(n606), .Z(n607) );
  NAND2_X1 U665 ( .A1(n700), .A2(n607), .ZN(n611) );
  NOR2_X1 U666 ( .A1(n599), .A2(n608), .ZN(n609) );
  XOR2_X1 U667 ( .A(KEYINPUT121), .B(n609), .Z(n610) );
  NOR2_X1 U668 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U669 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U670 ( .A(n614), .B(KEYINPUT122), .ZN(n615) );
  XOR2_X1 U671 ( .A(G143), .B(KEYINPUT117), .Z(n616) );
  XNOR2_X1 U672 ( .A(n617), .B(n616), .ZN(G45) );
  XNOR2_X1 U673 ( .A(n618), .B(G119), .ZN(G21) );
  XNOR2_X1 U674 ( .A(n619), .B(G101), .ZN(G3) );
  XNOR2_X1 U675 ( .A(n620), .B(KEYINPUT2), .ZN(n622) );
  NOR2_X4 U676 ( .A1(n622), .A2(n621), .ZN(n669) );
  NAND2_X1 U677 ( .A1(n669), .A2(G210), .ZN(n627) );
  XNOR2_X1 U678 ( .A(KEYINPUT91), .B(KEYINPUT54), .ZN(n623) );
  XNOR2_X1 U679 ( .A(n623), .B(KEYINPUT55), .ZN(n624) );
  XNOR2_X1 U680 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U681 ( .A(n627), .B(n626), .ZN(n629) );
  INV_X1 U682 ( .A(G952), .ZN(n628) );
  NOR2_X1 U683 ( .A1(n629), .A2(n678), .ZN(n631) );
  XOR2_X1 U684 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n630) );
  XNOR2_X1 U685 ( .A(n631), .B(n630), .ZN(G51) );
  INV_X1 U686 ( .A(KEYINPUT123), .ZN(n636) );
  NAND2_X1 U687 ( .A1(n669), .A2(G478), .ZN(n633) );
  XNOR2_X1 U688 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X1 U689 ( .A1(n634), .A2(n678), .ZN(n635) );
  XNOR2_X1 U690 ( .A(n636), .B(n635), .ZN(G63) );
  NAND2_X1 U691 ( .A1(n669), .A2(G472), .ZN(n640) );
  XOR2_X1 U692 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n637) );
  XNOR2_X1 U693 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U694 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X1 U695 ( .A1(n641), .A2(n678), .ZN(n643) );
  INV_X1 U696 ( .A(KEYINPUT63), .ZN(n642) );
  XNOR2_X1 U697 ( .A(n643), .B(n642), .ZN(G57) );
  XOR2_X1 U698 ( .A(G104), .B(KEYINPUT115), .Z(n646) );
  INV_X1 U699 ( .A(n644), .ZN(n657) );
  NAND2_X1 U700 ( .A1(n340), .A2(n657), .ZN(n645) );
  XNOR2_X1 U701 ( .A(n646), .B(n645), .ZN(G6) );
  XNOR2_X1 U702 ( .A(G107), .B(KEYINPUT27), .ZN(n651) );
  XOR2_X1 U703 ( .A(KEYINPUT116), .B(KEYINPUT26), .Z(n649) );
  INV_X1 U704 ( .A(n647), .ZN(n659) );
  NAND2_X1 U705 ( .A1(n340), .A2(n659), .ZN(n648) );
  XNOR2_X1 U706 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U707 ( .A(n651), .B(n650), .ZN(G9) );
  XNOR2_X1 U708 ( .A(G110), .B(n652), .ZN(G12) );
  XOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .Z(n654) );
  NAND2_X1 U710 ( .A1(n655), .A2(n659), .ZN(n653) );
  XNOR2_X1 U711 ( .A(n654), .B(n653), .ZN(G30) );
  NAND2_X1 U712 ( .A1(n655), .A2(n657), .ZN(n656) );
  XNOR2_X1 U713 ( .A(n656), .B(G146), .ZN(G48) );
  NAND2_X1 U714 ( .A1(n660), .A2(n657), .ZN(n658) );
  XNOR2_X1 U715 ( .A(n658), .B(G113), .ZN(G15) );
  NAND2_X1 U716 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U717 ( .A(n661), .B(G116), .ZN(G18) );
  XOR2_X1 U718 ( .A(G125), .B(KEYINPUT37), .Z(n662) );
  XNOR2_X1 U719 ( .A(n663), .B(n662), .ZN(G27) );
  NAND2_X1 U720 ( .A1(n669), .A2(G469), .ZN(n667) );
  XOR2_X1 U721 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n664) );
  NOR2_X1 U722 ( .A1(n668), .A2(n678), .ZN(G54) );
  NAND2_X1 U723 ( .A1(n669), .A2(G475), .ZN(n672) );
  XOR2_X1 U724 ( .A(n670), .B(KEYINPUT59), .Z(n671) );
  XNOR2_X1 U725 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U726 ( .A1(n673), .A2(n678), .ZN(n674) );
  XNOR2_X1 U727 ( .A(n674), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n669), .A2(G217), .ZN(n676) );
  XNOR2_X1 U729 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U730 ( .A1(n678), .A2(n677), .ZN(G66) );
  XNOR2_X1 U731 ( .A(n680), .B(n679), .ZN(n682) );
  NOR2_X1 U732 ( .A1(n700), .A2(G898), .ZN(n681) );
  NOR2_X1 U733 ( .A1(n682), .A2(n681), .ZN(n691) );
  NOR2_X1 U734 ( .A1(n683), .A2(G953), .ZN(n688) );
  INV_X1 U735 ( .A(G898), .ZN(n686) );
  NAND2_X1 U736 ( .A1(G953), .A2(G224), .ZN(n684) );
  XOR2_X1 U737 ( .A(KEYINPUT61), .B(n684), .Z(n685) );
  NOR2_X1 U738 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U739 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U740 ( .A(n689), .B(KEYINPUT124), .Z(n690) );
  XNOR2_X1 U741 ( .A(n691), .B(n690), .ZN(G69) );
  XOR2_X1 U742 ( .A(n693), .B(n692), .Z(n699) );
  XNOR2_X1 U743 ( .A(G227), .B(n699), .ZN(n694) );
  NAND2_X1 U744 ( .A1(n694), .A2(G900), .ZN(n695) );
  XOR2_X1 U745 ( .A(KEYINPUT125), .B(n695), .Z(n696) );
  NAND2_X1 U746 ( .A1(G953), .A2(n696), .ZN(n697) );
  XNOR2_X1 U747 ( .A(n697), .B(KEYINPUT126), .ZN(n703) );
  XNOR2_X1 U748 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U749 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U750 ( .A1(n703), .A2(n702), .ZN(G72) );
  XOR2_X1 U751 ( .A(G134), .B(n704), .Z(G36) );
  XOR2_X1 U752 ( .A(n705), .B(G137), .Z(G39) );
  XNOR2_X1 U753 ( .A(n706), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U754 ( .A(G140), .B(n707), .ZN(n708) );
  XNOR2_X1 U755 ( .A(n708), .B(KEYINPUT118), .ZN(G42) );
  XOR2_X1 U756 ( .A(G131), .B(n709), .Z(G33) );
endmodule

