//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  OAI211_X1 g003(.A(new_n188), .B(G146), .C1(new_n189), .C2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT82), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n195), .A3(new_n192), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT67), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n188), .A2(G146), .ZN(new_n201));
  AND4_X1   g015(.A1(KEYINPUT67), .A2(new_n198), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n194), .B(new_n196), .C1(new_n199), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(G107), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT10), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n205), .A2(new_n208), .A3(new_n210), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT81), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n223), .A3(G101), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n224), .A4(new_n211), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n200), .A2(new_n201), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n197), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n231), .A3(G101), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT65), .B(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n237), .A3(new_n239), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n193), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n199), .B2(new_n202), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n219), .A2(new_n234), .A3(new_n246), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G227), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT80), .ZN(new_n254));
  XNOR2_X1  g068(.A(G110), .B(G140), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n254), .B(new_n255), .Z(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n190), .A2(new_n195), .A3(new_n192), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n195), .B1(new_n190), .B2(new_n192), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n197), .A2(KEYINPUT67), .A3(new_n198), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n215), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n249), .B1(new_n266), .B2(KEYINPUT10), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n230), .A2(new_n232), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n220), .A2(new_n223), .A3(G101), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n211), .A2(KEYINPUT4), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(new_n222), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n245), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n257), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n251), .B1(new_n250), .B2(new_n256), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n248), .A2(new_n216), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT12), .B(new_n245), .C1(new_n277), .C2(new_n266), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT83), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n193), .B1(new_n263), .B2(new_n264), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n215), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n217), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT12), .A4(new_n245), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n245), .B1(new_n277), .B2(new_n266), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n256), .B1(new_n288), .B2(new_n250), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n276), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G469), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n250), .A2(new_n256), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n256), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n280), .A2(new_n218), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n217), .A2(new_n218), .B1(new_n295), .B2(new_n216), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n246), .B1(new_n296), .B2(new_n234), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n267), .A2(new_n272), .A3(new_n245), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT85), .B(G469), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT86), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n273), .A2(new_n250), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n288), .A2(new_n292), .B1(new_n304), .B2(new_n294), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n306));
  NOR4_X1   g120(.A1(new_n305), .A2(new_n306), .A3(G902), .A4(new_n301), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n291), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n312));
  NOR2_X1   g126(.A1(G475), .A2(G902), .ZN(new_n313));
  XNOR2_X1  g127(.A(G125), .B(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  OR3_X1    g130(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(G146), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(G146), .B1(new_n315), .B2(new_n317), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G237), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  OAI211_X1 g139(.A(G214), .B(new_n252), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n188), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(G237), .ZN(new_n329));
  AOI21_X1  g143(.A(G953), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G143), .A3(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT65), .B(G131), .Z(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n327), .A2(new_n243), .A3(new_n331), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n243), .B1(new_n327), .B2(new_n331), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT93), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT17), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n338), .B2(KEYINPUT17), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n321), .B(new_n337), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G113), .B(G122), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n204), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n314), .A2(new_n191), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT77), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n191), .B2(new_n314), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n332), .A2(KEYINPUT18), .A3(G131), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT18), .A2(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n327), .A2(new_n331), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n342), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n334), .A2(new_n336), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n334), .A2(KEYINPUT92), .A3(new_n336), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n314), .B(KEYINPUT19), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n319), .B1(new_n191), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n344), .B1(new_n359), .B2(new_n351), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n312), .B(new_n313), .C1(new_n352), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n313), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n358), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT92), .B1(new_n334), .B2(new_n336), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n351), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n344), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n342), .A2(new_n344), .A3(new_n351), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT94), .A3(new_n312), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n313), .B1(new_n352), .B2(new_n360), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT20), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n363), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n188), .A2(G128), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n188), .A2(G128), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n377), .A2(new_n378), .A3(G134), .ZN(new_n379));
  XNOR2_X1  g193(.A(G116), .B(G122), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n380), .A2(new_n207), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n207), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n376), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n385), .A2(KEYINPUT95), .B1(KEYINPUT13), .B2(new_n377), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(KEYINPUT95), .B2(new_n385), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n383), .B1(new_n387), .B2(G134), .ZN(new_n388));
  INV_X1    g202(.A(G116), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT14), .A3(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(new_n380), .ZN(new_n393));
  OAI21_X1  g207(.A(G134), .B1(new_n377), .B2(new_n378), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n381), .B(new_n393), .C1(new_n379), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n309), .A2(new_n396), .A3(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OR3_X1    g212(.A1(new_n388), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n388), .B2(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n187), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G478), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(G478), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n187), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n344), .B1(new_n342), .B2(new_n351), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n187), .B1(new_n352), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G475), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n375), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n311), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n414));
  INV_X1    g228(.A(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G128), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n415), .A2(G128), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(KEYINPUT23), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G110), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(KEYINPUT74), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n415), .A3(G128), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n421), .B(new_n423), .C1(new_n415), .C2(G128), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT24), .B(G110), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n321), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n346), .A2(new_n318), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n425), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT76), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n425), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT75), .B1(new_n419), .B2(G110), .ZN(new_n434));
  OR3_X1    g248(.A1(new_n419), .A2(KEYINPUT75), .A3(G110), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT78), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT22), .B(G137), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n428), .B2(new_n437), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n414), .B(new_n187), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(G217), .A2(G902), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n396), .B2(G234), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT73), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n442), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n414), .B1(new_n451), .B2(new_n187), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n413), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n443), .A2(new_n444), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT25), .B1(new_n454), .B2(G902), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT79), .A3(new_n448), .A4(new_n445), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n448), .A2(G902), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n236), .A2(G137), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n238), .A2(G134), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n241), .B2(new_n333), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n463), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n248), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT64), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n229), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n227), .B(KEYINPUT64), .C1(new_n197), .C2(new_n228), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n245), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G116), .B(G119), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT2), .B(G113), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(KEYINPUT2), .B(G113), .Z(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n464), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n248), .A2(new_n483), .B1(new_n245), .B2(new_n230), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT68), .B1(new_n484), .B2(KEYINPUT30), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n464), .B1(new_n265), .B2(new_n247), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n229), .B1(new_n244), .B2(new_n242), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n488));
  NOR4_X1   g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n474), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n475), .B(new_n482), .C1(new_n485), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n330), .A2(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n482), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n484), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT31), .ZN(new_n500));
  INV_X1    g314(.A(new_n496), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n473), .A2(new_n482), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n484), .A2(KEYINPUT28), .A3(new_n497), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT31), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n490), .A2(new_n508), .A3(new_n496), .A4(new_n498), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(G472), .A2(G902), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n460), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n460), .A3(new_n511), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n501), .B2(new_n506), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n490), .A2(new_n498), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n501), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n498), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT72), .B(new_n482), .C1(new_n486), .C2(new_n487), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(KEYINPUT28), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n503), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n496), .A2(KEYINPUT29), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n187), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G472), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n459), .B1(new_n515), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G210), .B1(G237), .B2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n280), .A2(new_n316), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n229), .A2(G125), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n252), .A2(G224), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n481), .A2(new_n211), .A3(new_n214), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT5), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n415), .A3(G116), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT87), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n541), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n542), .A2(new_n543), .A3(G113), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G122), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n223), .B1(new_n220), .B2(G101), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n269), .A2(new_n548), .A3(new_n270), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n482), .A2(new_n232), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT6), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(new_n547), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n554), .A2(new_n552), .A3(KEYINPUT6), .A4(new_n555), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n536), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n547), .B(KEYINPUT8), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n543), .B(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n542), .A2(G113), .A3(new_n544), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n537), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n216), .B1(new_n481), .B2(new_n545), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n532), .A2(KEYINPUT7), .A3(new_n533), .A4(new_n535), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n551), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n532), .A2(KEYINPUT90), .B1(G125), .B2(new_n229), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n570), .B1(KEYINPUT7), .B2(new_n535), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n187), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n531), .B1(new_n559), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n552), .A2(KEYINPUT6), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n482), .A2(new_n232), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(new_n225), .B1(new_n538), .B2(new_n545), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n576), .B2(new_n547), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n547), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n558), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n536), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n566), .A2(new_n551), .A3(new_n567), .ZN(new_n582));
  INV_X1    g396(.A(new_n571), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n584), .A3(new_n530), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n573), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT91), .B(new_n531), .C1(new_n559), .C2(new_n572), .ZN(new_n588));
  INV_X1    g402(.A(G952), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(G953), .ZN(new_n590));
  NAND2_X1  g404(.A1(G234), .A2(G237), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT21), .B(G898), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(G902), .A3(G953), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT96), .ZN(new_n597));
  OAI21_X1  g411(.A(G214), .B1(G237), .B2(G902), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n587), .A2(new_n588), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n412), .A2(new_n529), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT97), .B(G101), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G3));
  AND3_X1   g417(.A1(new_n453), .A2(new_n456), .A3(new_n458), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n510), .A2(new_n187), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n605), .A2(G472), .B1(new_n511), .B2(new_n510), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n604), .A2(new_n606), .A3(new_n308), .A4(new_n310), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT98), .ZN(new_n608));
  INV_X1    g422(.A(new_n310), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n279), .A2(new_n284), .A3(new_n287), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n250), .A2(new_n256), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n299), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n187), .A3(new_n302), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n306), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n300), .A2(KEYINPUT86), .A3(new_n302), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n609), .B1(new_n616), .B2(new_n291), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n604), .A4(new_n606), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n399), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n401), .A2(new_n622), .A3(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n399), .B(new_n400), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(G478), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(G478), .A2(G902), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n626), .B(new_n627), .C1(G478), .C2(new_n402), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n375), .B2(new_n410), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n573), .A2(new_n585), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n631), .B2(new_n598), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n598), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n573), .B2(new_n585), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n630), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n629), .A2(new_n633), .A3(new_n597), .A4(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n620), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G104), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n410), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n371), .A2(new_n645), .A3(new_n312), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n409), .A2(KEYINPUT103), .A3(G475), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n374), .A2(KEYINPUT102), .A3(new_n361), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n648), .A2(new_n649), .A3(new_n407), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT99), .B(new_n634), .C1(new_n573), .C2(new_n585), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n632), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n652), .A3(new_n597), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n620), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(new_n606), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n428), .A2(new_n437), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n441), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n457), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n453), .A2(new_n456), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n412), .A2(new_n665), .A3(new_n600), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NOR3_X1   g482(.A1(new_n311), .A2(new_n651), .A3(new_n632), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n510), .A2(new_n460), .A3(new_n511), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n528), .B1(new_n670), .B2(new_n512), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n663), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n595), .A2(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n592), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n650), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT104), .B(G128), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G30));
  XNOR2_X1  g493(.A(new_n675), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n617), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT40), .Z(new_n682));
  AOI21_X1  g496(.A(new_n501), .B1(new_n498), .B2(new_n490), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n522), .A2(new_n523), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n187), .B1(new_n684), .B2(new_n496), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n670), .B2(new_n512), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n587), .A2(new_n588), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n407), .B1(new_n375), .B2(new_n410), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n664), .A2(new_n692), .A3(new_n598), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n682), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND2_X1  g510(.A1(new_n629), .A2(new_n675), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n673), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT106), .B(G146), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G48));
  NAND2_X1  g514(.A1(new_n671), .A2(new_n604), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n637), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n305), .B2(G902), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n310), .B(new_n703), .C1(new_n303), .C2(new_n307), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n616), .A2(new_n706), .A3(new_n310), .A4(new_n703), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n705), .A2(new_n707), .A3(KEYINPUT108), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n702), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NOR2_X1   g528(.A1(new_n653), .A2(new_n701), .ZN(new_n715));
  AND4_X1   g529(.A1(KEYINPUT109), .A2(new_n715), .A3(new_n711), .A4(new_n710), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n705), .A2(new_n707), .A3(KEYINPUT108), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n705), .B2(new_n707), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT109), .B1(new_n719), .B2(new_n715), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n389), .ZN(G18));
  NAND3_X1  g536(.A1(new_n705), .A2(new_n652), .A3(new_n707), .ZN(new_n723));
  INV_X1    g537(.A(new_n411), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n671), .A3(new_n597), .A4(new_n663), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n415), .ZN(G21));
  NAND3_X1  g541(.A1(new_n605), .A2(KEYINPUT111), .A3(G472), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n525), .A2(new_n501), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n500), .A2(new_n729), .A3(new_n509), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT110), .B1(new_n730), .B2(new_n511), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(KEYINPUT110), .A3(new_n511), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT111), .B1(new_n605), .B2(G472), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n459), .A3(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n652), .A2(new_n597), .A3(new_n692), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n710), .A2(new_n736), .A3(new_n737), .A4(new_n711), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  AND3_X1   g553(.A1(new_n705), .A2(new_n652), .A3(new_n707), .ZN(new_n740));
  INV_X1    g554(.A(new_n733), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n731), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n605), .A2(G472), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n745), .A3(new_n663), .A4(new_n728), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n697), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n740), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n634), .B1(new_n587), .B2(new_n588), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n617), .A2(new_n671), .A3(new_n604), .A4(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n753), .B2(new_n697), .ZN(new_n754));
  INV_X1    g568(.A(new_n752), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n311), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n529), .A2(new_n756), .A3(new_n748), .A4(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  OAI21_X1  g573(.A(KEYINPUT112), .B1(new_n753), .B2(new_n676), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n761));
  INV_X1    g575(.A(new_n675), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n648), .A2(new_n649), .A3(new_n407), .A4(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n756), .A2(new_n529), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n276), .A2(new_n289), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n276), .B2(new_n289), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(G469), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(G469), .A2(G902), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n614), .B2(new_n615), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n771), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n609), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n680), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n375), .A2(new_n410), .ZN(new_n777));
  INV_X1    g591(.A(new_n628), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n375), .A2(new_n410), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n781), .A2(KEYINPUT43), .A3(new_n628), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n658), .A3(new_n663), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n755), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n776), .B(new_n785), .C1(new_n784), .C2(new_n783), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NOR4_X1   g601(.A1(new_n697), .A2(new_n671), .A3(new_n755), .A4(new_n604), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n790), .B(new_n609), .C1(new_n773), .C2(new_n774), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n589), .A2(new_n252), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n708), .A2(new_n755), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n687), .B(KEYINPUT105), .ZN(new_n797));
  INV_X1    g611(.A(new_n592), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n604), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n781), .A3(new_n778), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n780), .A2(new_n798), .A3(new_n782), .ZN(new_n802));
  INV_X1    g616(.A(new_n736), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n691), .A2(new_n634), .ZN(new_n805));
  INV_X1    g619(.A(new_n708), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n801), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n802), .A2(new_n803), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(KEYINPUT50), .A3(new_n806), .A4(new_n805), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n800), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n705), .A2(new_n707), .A3(new_n752), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n802), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n802), .B2(new_n813), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n747), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n816), .B2(new_n747), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n795), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n747), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT119), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n811), .A3(KEYINPUT120), .A4(new_n818), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n616), .A2(new_n609), .A3(new_n703), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n804), .A2(new_n755), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n821), .A2(new_n824), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n629), .ZN(new_n833));
  OAI221_X1 g647(.A(new_n590), .B1(new_n799), .B2(new_n833), .C1(new_n804), .C2(new_n723), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT121), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT48), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n816), .B(new_n529), .C1(KEYINPUT122), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(KEYINPUT122), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n826), .A2(KEYINPUT116), .A3(new_n827), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n789), .B2(new_n791), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n844), .A3(new_n828), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n845), .A2(new_n846), .A3(new_n830), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n823), .A2(new_n811), .A3(new_n818), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n845), .B2(new_n830), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n832), .B(new_n841), .C1(new_n850), .C2(KEYINPUT51), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n819), .A2(new_n820), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n830), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n825), .B1(new_n857), .B2(new_n847), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(KEYINPUT123), .A3(new_n832), .A4(new_n841), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n652), .A2(new_n692), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n311), .A2(new_n663), .A3(new_n762), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n689), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n669), .B(new_n672), .C1(new_n763), .C2(new_n748), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n749), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT52), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n864), .A2(new_n749), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n867), .A2(KEYINPUT115), .A3(new_n869), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n726), .B1(new_n719), .B2(new_n702), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n738), .B(new_n876), .C1(new_n716), .C2(new_n720), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n629), .A2(new_n600), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT113), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n629), .A2(new_n600), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n608), .A2(new_n619), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n412), .B(new_n600), .C1(new_n529), .C2(new_n665), .ZN(new_n883));
  INV_X1    g697(.A(new_n407), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n777), .A2(new_n600), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n608), .A2(new_n619), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n754), .A2(new_n757), .B1(new_n760), .B2(new_n764), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n407), .A2(new_n675), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n648), .A2(new_n649), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n671), .A3(new_n663), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n746), .B2(new_n697), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n756), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n875), .B1(new_n877), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n723), .A2(new_n725), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n738), .A2(new_n712), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n719), .A2(new_n715), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT109), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n719), .A2(KEYINPUT109), .A3(new_n715), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n758), .A2(new_n765), .A3(new_n893), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT114), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n895), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n874), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n870), .B1(new_n895), .B2(new_n906), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n908), .B(KEYINPUT54), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n872), .A2(new_n873), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n877), .A2(new_n894), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n914), .B(new_n915), .C1(new_n910), .C2(KEYINPUT53), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n794), .B1(new_n860), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n616), .A2(new_n703), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT49), .Z(new_n920));
  NOR4_X1   g734(.A1(new_n779), .A2(new_n459), .A3(new_n634), .A4(new_n609), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n921), .A3(new_n797), .A4(new_n691), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n922), .ZN(G75));
  INV_X1    g737(.A(new_n870), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n877), .A2(new_n894), .A3(new_n875), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT114), .B1(new_n902), .B2(new_n905), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n909), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n914), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n579), .B(new_n580), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n252), .A2(G952), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G51));
  NOR2_X1   g752(.A1(new_n910), .A2(KEYINPUT53), .ZN(new_n939));
  INV_X1    g753(.A(new_n914), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT54), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n916), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n771), .B(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT57), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n612), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n939), .A2(new_n940), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n947), .A2(new_n187), .A3(new_n770), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n937), .B1(new_n946), .B2(new_n948), .ZN(G54));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n187), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n369), .A2(new_n370), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n937), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n950), .A2(KEYINPUT58), .A3(G475), .A4(new_n952), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(G60));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n623), .A2(new_n625), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n627), .B(KEYINPUT59), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n915), .B1(new_n928), .B2(new_n914), .ZN(new_n964));
  INV_X1    g778(.A(new_n916), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n955), .ZN(new_n967));
  INV_X1    g781(.A(new_n962), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n960), .B1(new_n917), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n958), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n917), .A2(new_n968), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n961), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n937), .B1(new_n942), .B2(new_n963), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(G63));
  XNOR2_X1  g789(.A(new_n446), .B(KEYINPUT60), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n454), .B1(new_n947), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n929), .A2(new_n661), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n955), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G66));
  AOI21_X1  g796(.A(new_n252), .B1(new_n594), .B2(G224), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n877), .A2(new_n904), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n985), .B2(new_n252), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n557), .B(new_n558), .C1(G898), .C2(new_n252), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(G69));
  NOR2_X1   g802(.A1(new_n485), .A2(new_n489), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n474), .B2(new_n473), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n357), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n629), .B1(new_n884), .B2(new_n777), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n992), .A2(new_n681), .A3(new_n701), .A4(new_n755), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n786), .A2(new_n792), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n749), .A2(new_n865), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n695), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n993), .B(new_n994), .C1(KEYINPUT62), .C2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n991), .B1(new_n999), .B2(new_n252), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n776), .A2(new_n529), .A3(new_n862), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n995), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(new_n786), .A3(new_n792), .A4(new_n888), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(G953), .ZN(new_n1004));
  INV_X1    g818(.A(G900), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n991), .B1(new_n1005), .B2(new_n252), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n252), .B1(G227), .B2(G900), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n1003), .B2(new_n985), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n518), .A2(new_n496), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n937), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n997), .A2(new_n984), .A3(new_n998), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1016), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n683), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g835(.A1(new_n927), .A2(KEYINPUT53), .B1(new_n907), .B2(new_n874), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1012), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1014), .A2(new_n683), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(G57));
endmodule


