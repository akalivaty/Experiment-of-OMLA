//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT91), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G137), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n193), .B2(G137), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n192), .A3(new_n197), .A4(new_n194), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(new_n199), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n200), .A2(new_n202), .B1(new_n203), .B2(G131), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT88), .B1(new_n205), .B2(G104), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G104), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G107), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n205), .A2(KEYINPUT3), .A3(G104), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT3), .B1(new_n205), .B2(G104), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT10), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT64), .B1(new_n220), .B2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT1), .B1(new_n220), .B2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(G143), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n230), .A2(new_n225), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n219), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n218), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n225), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .A3(new_n232), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n230), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(G128), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n212), .A2(new_n217), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n236), .B1(new_n245), .B2(KEYINPUT10), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(KEYINPUT0), .A3(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G101), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT0), .B(G128), .Z(new_n252));
  AND3_X1   g066(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT65), .B1(new_n226), .B2(new_n252), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n248), .B(new_n251), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT86), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n208), .B2(G107), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n205), .A2(KEYINPUT3), .A3(G104), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n213), .B1(new_n262), .B2(new_n214), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n257), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n260), .A2(new_n261), .B1(new_n208), .B2(G107), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n250), .B1(new_n265), .B2(new_n213), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n249), .A2(G101), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(KEYINPUT86), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n256), .A2(new_n269), .A3(KEYINPUT87), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT87), .B1(new_n256), .B2(new_n269), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n204), .B(new_n247), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G227), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(KEYINPUT90), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n203), .A2(G131), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n229), .A2(new_n234), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n218), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n245), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT90), .B1(new_n272), .B2(new_n277), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n190), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n272), .A2(new_n277), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT90), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n293), .A2(KEYINPUT91), .A3(new_n287), .A4(new_n278), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n247), .B1(new_n270), .B2(new_n271), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n295), .A2(new_n282), .ZN(new_n296));
  INV_X1    g110(.A(new_n272), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n276), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n290), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n287), .A2(new_n272), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n303), .A2(new_n277), .B1(new_n291), .B2(new_n296), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(new_n300), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n189), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G113), .B(G122), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(new_n208), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n312), .A2(KEYINPUT78), .A3(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT78), .B1(new_n312), .B2(G140), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n314), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G146), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G214), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(new_n220), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT18), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n197), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n326), .B(G143), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT18), .A3(G131), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n311), .A2(new_n323), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n315), .A2(G125), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n316), .A3(KEYINPUT81), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n333), .B2(new_n313), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n223), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT95), .A3(new_n322), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n310), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n321), .A2(KEYINPUT16), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n313), .A2(KEYINPUT16), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n223), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n327), .A2(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n330), .A2(new_n197), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT19), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n349), .A3(new_n337), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n321), .B2(new_n349), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n223), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(G475), .A2(G902), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT17), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n346), .A2(new_n347), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n356), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n342), .A2(new_n223), .A3(new_n343), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n344), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n359), .A2(new_n361), .B1(new_n340), .B2(new_n332), .ZN(new_n362));
  INV_X1    g176(.A(new_n310), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n354), .B(new_n355), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT20), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n359), .A2(new_n361), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n332), .A2(new_n340), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n310), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n354), .A4(new_n355), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n310), .A2(KEYINPUT96), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n301), .B1(new_n368), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g189(.A(G475), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n232), .A2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n232), .A2(G143), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(KEYINPUT13), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n193), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n220), .A2(G128), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT97), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n382), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n383), .A2(new_n379), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n193), .ZN(new_n388));
  XNOR2_X1  g202(.A(G116), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n205), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n387), .B(new_n193), .ZN(new_n392));
  INV_X1    g206(.A(G116), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT14), .A3(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n389), .ZN(new_n395));
  OAI211_X1 g209(.A(G107), .B(new_n394), .C1(new_n395), .C2(KEYINPUT14), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n392), .B(new_n396), .C1(G107), .C2(new_n395), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n187), .A2(new_n399), .A3(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n391), .B2(new_n397), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n301), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT15), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n404), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT21), .B(G898), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT98), .ZN(new_n410));
  NAND2_X1  g224(.A1(G234), .A2(G237), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n411), .A2(G902), .A3(G953), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n411), .A2(G952), .A3(new_n325), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT99), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n377), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT8), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT2), .B(G113), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G116), .B(G119), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n425));
  INV_X1    g239(.A(G119), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G116), .ZN(new_n427));
  INV_X1    g241(.A(new_n423), .ZN(new_n428));
  OAI211_X1 g242(.A(G113), .B(new_n427), .C1(new_n428), .C2(new_n425), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n424), .A2(new_n429), .A3(new_n217), .A4(new_n212), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n429), .A2(new_n424), .B1(new_n212), .B2(new_n217), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n420), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n283), .A2(G125), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(G125), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n325), .A2(G224), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(KEYINPUT7), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n437), .B2(KEYINPUT7), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n432), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n428), .A2(new_n421), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n424), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n251), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n264), .B2(new_n268), .ZN(new_n444));
  INV_X1    g258(.A(new_n419), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n445), .A3(new_n430), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(KEYINPUT7), .A3(new_n436), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n448), .A2(new_n449), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n430), .ZN(new_n453));
  INV_X1    g267(.A(new_n269), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n419), .B(new_n453), .C1(new_n454), .C2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n445), .B1(new_n444), .B2(new_n430), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT6), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n435), .B(new_n436), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n459), .B(new_n445), .C1(new_n444), .C2(new_n430), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n461), .A3(new_n301), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n452), .A2(new_n461), .A3(new_n301), .A4(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G214), .B1(G237), .B2(G902), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT92), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n418), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n308), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G472), .A2(G902), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT26), .B(G101), .Z(new_n475));
  NAND3_X1  g289(.A1(new_n324), .A2(new_n325), .A3(G210), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n191), .A2(G134), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n197), .B1(new_n480), .B2(new_n194), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n229), .B2(new_n234), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n200), .A2(new_n202), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n434), .B2(new_n204), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n442), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n231), .A2(KEYINPUT0), .A3(G128), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n226), .A2(new_n252), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n252), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n282), .ZN(new_n493));
  INV_X1    g307(.A(new_n442), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n484), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n479), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT67), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n434), .A2(new_n204), .ZN(new_n504));
  INV_X1    g318(.A(new_n481), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n283), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n201), .B(new_n196), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT30), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n442), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT30), .B1(new_n493), .B2(new_n484), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n482), .B2(new_n483), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n494), .B1(new_n493), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n485), .A2(new_n512), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT67), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n495), .A2(new_n479), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT31), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n521), .B(new_n518), .C1(new_n511), .C2(new_n516), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n502), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT67), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT67), .B1(new_n514), .B2(new_n515), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n521), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(KEYINPUT31), .A3(new_n519), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT70), .A3(new_n502), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n474), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT71), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n534));
  INV_X1    g348(.A(G472), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n517), .A2(new_n495), .ZN(new_n536));
  INV_X1    g350(.A(new_n479), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n496), .A2(new_n497), .B1(new_n499), .B2(new_n495), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT29), .B1(new_n539), .B2(new_n479), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n496), .A2(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT72), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n495), .A2(KEYINPUT73), .A3(new_n499), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT73), .B1(new_n495), .B2(new_n499), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT72), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n496), .A2(new_n547), .A3(KEYINPUT28), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n479), .A2(KEYINPUT29), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n535), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT70), .B1(new_n531), .B2(new_n502), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n524), .B(new_n501), .C1(new_n529), .C2(new_n530), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n473), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT71), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n534), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT80), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G110), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n426), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n232), .A2(G119), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT74), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT74), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT79), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n568));
  AOI22_X1  g382(.A1(KEYINPUT76), .A2(new_n568), .B1(new_n232), .B2(G119), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(KEYINPUT76), .B2(new_n568), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n570), .A2(new_n563), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n567), .B1(new_n575), .B2(G110), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n561), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n574), .A2(new_n573), .ZN(new_n582));
  INV_X1    g396(.A(G110), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n563), .A4(new_n570), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT80), .A3(new_n579), .A4(new_n567), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n345), .A3(new_n339), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n575), .A2(G110), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n565), .A2(new_n566), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(new_n562), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n361), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT82), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n587), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n345), .A2(new_n339), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n581), .B2(new_n585), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n600), .B2(new_n591), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT25), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n399), .B1(G234), .B2(new_n301), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT83), .B1(new_n605), .B2(KEYINPUT25), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n602), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(G902), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n597), .A2(new_n601), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n608), .A2(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n472), .A2(new_n560), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NAND2_X1  g432(.A1(new_n525), .A2(new_n532), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n535), .B1(new_n619), .B2(new_n301), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n533), .ZN(new_n621));
  INV_X1    g435(.A(new_n467), .ZN(new_n622));
  INV_X1    g436(.A(new_n468), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n621), .A2(new_n616), .A3(new_n308), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n405), .A2(new_n301), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n627), .B1(new_n404), .B2(G478), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n398), .B(new_n401), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n631), .B2(G478), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n372), .A2(new_n376), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n417), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  XNOR2_X1  g454(.A(new_n404), .B(new_n406), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n372), .A2(new_n376), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n417), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n625), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n587), .A2(new_n592), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n614), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT25), .B1(new_n604), .B2(new_n605), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(new_n611), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n472), .A2(new_n621), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT101), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G12));
  NAND2_X1  g472(.A1(new_n624), .A2(new_n654), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n414), .B1(new_n412), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n643), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n560), .A2(new_n308), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XOR2_X1   g480(.A(new_n661), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n308), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n536), .A2(new_n479), .ZN(new_n671));
  INV_X1    g485(.A(new_n496), .ZN(new_n672));
  AOI21_X1  g486(.A(G902), .B1(new_n672), .B2(new_n537), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n535), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n534), .A2(new_n675), .A3(new_n559), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT38), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n467), .B(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n408), .B1(new_n372), .B2(new_n376), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n468), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n678), .A2(new_n654), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n669), .A2(new_n670), .A3(new_n676), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND3_X1  g497(.A1(new_n632), .A2(new_n633), .A3(new_n662), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n659), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n560), .A2(new_n308), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND2_X1  g501(.A1(new_n299), .A2(new_n301), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n188), .A2(new_n689), .A3(new_n302), .A4(new_n624), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n560), .A2(new_n690), .A3(new_n616), .A4(new_n636), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NOR2_X1   g507(.A1(new_n642), .A2(new_n635), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n560), .A2(new_n690), .A3(new_n616), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NAND2_X1  g510(.A1(new_n689), .A2(new_n302), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n189), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n659), .A2(new_n418), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n560), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n529), .A2(new_n530), .B1(new_n549), .B2(new_n537), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n473), .B(KEYINPUT102), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n549), .A2(new_n537), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n531), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n704), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(KEYINPUT103), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n620), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n467), .A2(new_n679), .A3(new_n468), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n635), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n698), .A2(new_n616), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  INV_X1    g529(.A(new_n654), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n620), .A2(new_n716), .A3(new_n710), .ZN(new_n717));
  INV_X1    g531(.A(new_n684), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n690), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NOR2_X1   g534(.A1(new_n556), .A2(new_n558), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT105), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n552), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n556), .A2(new_n558), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT104), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n308), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n616), .A3(new_n718), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n560), .A2(new_n616), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n308), .A2(new_n731), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n733), .A2(KEYINPUT42), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  INV_X1    g553(.A(new_n663), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n732), .A2(new_n560), .A3(new_n616), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(new_n731), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n377), .A2(new_n632), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT43), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n621), .A2(new_n745), .A3(new_n716), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n743), .B1(new_n746), .B2(KEYINPUT44), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(KEYINPUT44), .B2(new_n746), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n304), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n300), .B1(new_n304), .B2(new_n749), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n306), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n302), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT107), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n756), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n302), .A4(new_n754), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n188), .A3(new_n667), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n748), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n191), .ZN(G39));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n188), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n762), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n560), .A2(new_n616), .A3(new_n743), .A4(new_n684), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  NOR2_X1   g587(.A1(new_n697), .A2(KEYINPUT49), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT108), .ZN(new_n775));
  INV_X1    g589(.A(new_n676), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n697), .A2(KEYINPUT49), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n188), .A2(new_n377), .A3(new_n469), .A4(new_n632), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n678), .A2(new_n616), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n665), .A2(new_n719), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n652), .B(new_n662), .C1(new_n653), .C2(new_n611), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n712), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n308), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n676), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n686), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n781), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n665), .A2(new_n686), .A3(new_n719), .A4(new_n786), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n782), .A2(new_n787), .A3(new_n781), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n716), .A2(new_n633), .A3(new_n641), .A4(new_n661), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n560), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n717), .A2(new_n718), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n735), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n560), .A2(new_n732), .A3(new_n616), .A4(new_n740), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n560), .A2(new_n798), .B1(new_n717), .B2(new_n718), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT110), .B(new_n741), .C1(new_n804), .C2(new_n735), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n691), .A2(new_n695), .A3(new_n700), .A4(new_n714), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n644), .B2(new_n470), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n694), .A2(KEYINPUT109), .A3(new_n467), .A4(new_n469), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n809), .B(new_n810), .C1(new_n470), .C2(new_n637), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n616), .A3(new_n308), .A4(new_n621), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n617), .A2(new_n812), .A3(new_n655), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n806), .A2(new_n738), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT53), .B1(new_n796), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n807), .B(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n733), .A2(KEYINPUT42), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n736), .A2(new_n737), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n788), .A2(new_n790), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n806), .A2(new_n818), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n816), .A2(new_n825), .A3(KEYINPUT54), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n678), .A2(new_n623), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n698), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n698), .A2(KEYINPUT113), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n745), .A2(new_n415), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n616), .A3(new_n711), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n835), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT114), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT50), .B1(new_n832), .B2(new_n835), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n837), .B(new_n834), .C1(new_n830), .C2(new_n831), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n698), .A2(new_n414), .A3(new_n731), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n745), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n717), .ZN(new_n848));
  INV_X1    g662(.A(new_n846), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n616), .A3(new_n776), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n632), .A2(new_n633), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n697), .A2(new_n188), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n768), .A2(new_n769), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n834), .A2(new_n743), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT51), .B1(new_n845), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  INV_X1    g673(.A(new_n852), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n838), .B2(new_n839), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(G952), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n864), .B(G953), .C1(new_n835), .C2(new_n690), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n634), .B2(new_n850), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n729), .A2(new_n616), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n847), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(KEYINPUT48), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(KEYINPUT48), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n858), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n815), .A2(new_n819), .A3(new_n824), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n806), .A2(new_n738), .A3(new_n814), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n791), .B2(new_n795), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n874), .B(KEYINPUT54), .C1(new_n876), .C2(new_n819), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n826), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n864), .A2(new_n325), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n780), .B1(new_n880), .B2(new_n882), .ZN(G75));
  NAND2_X1  g697(.A1(new_n864), .A2(G953), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT116), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n818), .A2(new_n823), .A3(new_n824), .A4(new_n806), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n876), .B2(KEYINPUT53), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(G210), .A3(G902), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n457), .A2(new_n460), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n458), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n894), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n886), .B1(new_n895), .B2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(new_n306), .B(KEYINPUT57), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n299), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n888), .A2(G902), .A3(new_n750), .A4(new_n751), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n886), .B1(new_n902), .B2(new_n903), .ZN(G54));
  NAND2_X1  g718(.A1(KEYINPUT58), .A2(G475), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT117), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n888), .A2(G902), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n369), .A2(new_n354), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n907), .A2(new_n909), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n886), .ZN(G60));
  NOR2_X1   g726(.A1(new_n899), .A2(new_n900), .ZN(new_n913));
  INV_X1    g727(.A(new_n631), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n627), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n885), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n826), .A2(new_n877), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n919), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT60), .Z(new_n923));
  OAI211_X1 g737(.A(new_n651), .B(new_n923), .C1(new_n816), .C2(new_n825), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT119), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n888), .A2(new_n926), .A3(new_n651), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n888), .A2(new_n923), .ZN(new_n929));
  INV_X1    g743(.A(new_n615), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n886), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(G66));
  INV_X1    g749(.A(G224), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n410), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n814), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n892), .B1(G898), .B2(new_n325), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  NAND2_X1  g754(.A1(new_n782), .A2(new_n686), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n682), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT62), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n634), .A2(new_n642), .ZN(new_n945));
  NOR4_X1   g759(.A1(new_n734), .A2(new_n668), .A3(new_n743), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n764), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n942), .A2(new_n948), .A3(new_n682), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n944), .A2(new_n772), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n325), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n515), .B1(new_n504), .B2(new_n508), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n351), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT121), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n738), .A2(new_n741), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT125), .Z(new_n957));
  NAND3_X1  g771(.A1(new_n867), .A2(new_n624), .A3(new_n679), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n763), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n770), .B2(new_n771), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n764), .B2(new_n941), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n942), .B(KEYINPUT124), .C1(new_n763), .C2(new_n748), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n957), .A2(new_n960), .A3(new_n964), .A4(new_n325), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n953), .B1(G900), .B2(G953), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n274), .B2(new_n660), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT122), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n954), .A2(KEYINPUT121), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n955), .A2(new_n967), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n967), .A2(new_n954), .ZN(new_n973));
  INV_X1    g787(.A(new_n969), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT126), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n976), .B(new_n969), .C1(new_n967), .C2(new_n954), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n972), .B1(new_n975), .B2(new_n977), .ZN(G72));
  XNOR2_X1  g792(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n535), .A2(new_n301), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n814), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n950), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n479), .A3(new_n536), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n874), .B1(new_n876), .B2(new_n819), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n538), .A2(new_n528), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n981), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n984), .B(new_n885), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n957), .A2(new_n964), .A3(new_n960), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n981), .B1(new_n989), .B2(new_n982), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n536), .A2(new_n479), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G57));
endmodule


