

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;

  XNOR2_X1 U324 ( .A(n336), .B(n327), .ZN(n328) );
  XNOR2_X1 U325 ( .A(n427), .B(KEYINPUT37), .ZN(n428) );
  XOR2_X1 U326 ( .A(n333), .B(n332), .Z(n540) );
  AND2_X1 U327 ( .A1(n572), .A2(n582), .ZN(n472) );
  XNOR2_X1 U328 ( .A(n430), .B(KEYINPUT73), .ZN(n431) );
  INV_X1 U329 ( .A(G176GAT), .ZN(n325) );
  XNOR2_X1 U330 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U331 ( .A(n483), .B(KEYINPUT48), .ZN(n534) );
  XNOR2_X1 U332 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U333 ( .A(n440), .B(n439), .ZN(n441) );
  INV_X1 U334 ( .A(n534), .ZN(n536) );
  INV_X1 U335 ( .A(KEYINPUT108), .ZN(n427) );
  XNOR2_X1 U336 ( .A(n442), .B(n441), .ZN(n448) );
  XNOR2_X1 U337 ( .A(n335), .B(KEYINPUT99), .ZN(n577) );
  NOR2_X1 U338 ( .A1(n383), .A2(n382), .ZN(n495) );
  INV_X1 U339 ( .A(n577), .ZN(n581) );
  XNOR2_X1 U340 ( .A(n429), .B(n428), .ZN(n524) );
  XOR2_X1 U341 ( .A(n587), .B(KEYINPUT41), .Z(n572) );
  INV_X1 U342 ( .A(G43GAT), .ZN(n469) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n491) );
  XNOR2_X1 U344 ( .A(n469), .B(KEYINPUT40), .ZN(n470) );
  XNOR2_X1 U345 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n471), .B(n470), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(G22GAT), .B(G155GAT), .Z(n397) );
  XOR2_X1 U348 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n293) );
  XNOR2_X1 U349 ( .A(KEYINPUT23), .B(G204GAT), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n397), .B(n294), .ZN(n296) );
  AND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n298) );
  INV_X1 U354 ( .A(KEYINPUT24), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n301) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(KEYINPUT79), .ZN(n299) );
  XOR2_X1 U357 ( .A(n299), .B(G162GAT), .Z(n422) );
  XOR2_X1 U358 ( .A(n422), .B(KEYINPUT93), .Z(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n304) );
  XOR2_X1 U360 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n303) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n350) );
  XOR2_X1 U363 ( .A(n304), .B(n350), .Z(n311) );
  XOR2_X1 U364 ( .A(KEYINPUT91), .B(G218GAT), .Z(n306) );
  XNOR2_X1 U365 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(n307), .ZN(n345) );
  XOR2_X1 U368 ( .A(G78GAT), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U369 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n435) );
  XOR2_X1 U371 ( .A(n345), .B(n435), .Z(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n485) );
  XOR2_X1 U373 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n313) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n333) );
  XOR2_X1 U376 ( .A(G190GAT), .B(G99GAT), .Z(n315) );
  XOR2_X1 U377 ( .A(G15GAT), .B(G127GAT), .Z(n398) );
  XOR2_X1 U378 ( .A(G113GAT), .B(KEYINPUT0), .Z(n347) );
  XNOR2_X1 U379 ( .A(n398), .B(n347), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U381 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XOR2_X1 U382 ( .A(n316), .B(n436), .Z(n331) );
  XOR2_X1 U383 ( .A(G183GAT), .B(KEYINPUT64), .Z(n318) );
  XNOR2_X1 U384 ( .A(KEYINPUT20), .B(KEYINPUT89), .ZN(n317) );
  XNOR2_X1 U385 ( .A(n318), .B(n317), .ZN(n329) );
  INV_X1 U386 ( .A(KEYINPUT17), .ZN(n319) );
  NAND2_X1 U387 ( .A1(n319), .A2(KEYINPUT19), .ZN(n322) );
  INV_X1 U388 ( .A(KEYINPUT19), .ZN(n320) );
  NAND2_X1 U389 ( .A1(n320), .A2(KEYINPUT17), .ZN(n321) );
  NAND2_X1 U390 ( .A1(n322), .A2(n321), .ZN(n324) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n323) );
  XNOR2_X1 U392 ( .A(n324), .B(n323), .ZN(n336) );
  NAND2_X1 U393 ( .A1(G227GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  NAND2_X1 U396 ( .A1(n485), .A2(n540), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n334), .B(KEYINPUT26), .ZN(n335) );
  XOR2_X1 U398 ( .A(KEYINPUT98), .B(n336), .Z(n338) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U401 ( .A(G8GAT), .B(G183GAT), .Z(n390) );
  XOR2_X1 U402 ( .A(n339), .B(n390), .Z(n344) );
  XOR2_X1 U403 ( .A(G92GAT), .B(G64GAT), .Z(n341) );
  XNOR2_X1 U404 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U406 ( .A(G176GAT), .B(n342), .Z(n446) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .Z(n408) );
  XNOR2_X1 U408 ( .A(n446), .B(n408), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n527) );
  XNOR2_X1 U411 ( .A(n527), .B(KEYINPUT27), .ZN(n379) );
  XOR2_X1 U412 ( .A(G134GAT), .B(KEYINPUT81), .Z(n409) );
  XOR2_X1 U413 ( .A(G85GAT), .B(n409), .Z(n349) );
  XNOR2_X1 U414 ( .A(n347), .B(G162GAT), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U416 ( .A(n350), .B(KEYINPUT96), .Z(n352) );
  NAND2_X1 U417 ( .A1(G225GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U419 ( .A(n354), .B(n353), .Z(n356) );
  XNOR2_X1 U420 ( .A(G29GAT), .B(G148GAT), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U422 ( .A(G57GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U423 ( .A(G120GAT), .B(G127GAT), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U425 ( .A(n360), .B(n359), .Z(n368) );
  XOR2_X1 U426 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n362) );
  XNOR2_X1 U427 ( .A(KEYINPUT97), .B(KEYINPUT95), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U429 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n364) );
  XNOR2_X1 U430 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n578) );
  INV_X1 U434 ( .A(n578), .ZN(n374) );
  NOR2_X1 U435 ( .A1(n379), .A2(n374), .ZN(n369) );
  NAND2_X1 U436 ( .A1(n577), .A2(n369), .ZN(n376) );
  XNOR2_X1 U437 ( .A(KEYINPUT25), .B(KEYINPUT100), .ZN(n372) );
  NOR2_X1 U438 ( .A1(n540), .A2(n527), .ZN(n370) );
  NOR2_X1 U439 ( .A1(n485), .A2(n370), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n373) );
  OR2_X1 U441 ( .A1(n374), .A2(n373), .ZN(n375) );
  NAND2_X1 U442 ( .A1(n376), .A2(n375), .ZN(n378) );
  INV_X1 U443 ( .A(KEYINPUT101), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U445 ( .A(n485), .B(KEYINPUT28), .Z(n538) );
  INV_X1 U446 ( .A(n538), .ZN(n381) );
  NOR2_X1 U447 ( .A1(n578), .A2(n379), .ZN(n535) );
  NAND2_X1 U448 ( .A1(n540), .A2(n535), .ZN(n380) );
  NOR2_X1 U449 ( .A1(n381), .A2(n380), .ZN(n382) );
  XOR2_X1 U450 ( .A(KEYINPUT86), .B(G64GAT), .Z(n385) );
  XNOR2_X1 U451 ( .A(G1GAT), .B(G71GAT), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n387) );
  XNOR2_X1 U454 ( .A(KEYINPUT14), .B(KEYINPUT83), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n402) );
  XOR2_X1 U457 ( .A(G57GAT), .B(KEYINPUT13), .Z(n433) );
  XOR2_X1 U458 ( .A(n390), .B(n433), .Z(n392) );
  XNOR2_X1 U459 ( .A(G211GAT), .B(G78GAT), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U461 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n394) );
  NAND2_X1 U462 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U463 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U464 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U467 ( .A(n402), .B(n401), .Z(n563) );
  INV_X1 U468 ( .A(n563), .ZN(n592) );
  NOR2_X1 U469 ( .A1(n495), .A2(n592), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n403), .B(KEYINPUT107), .ZN(n426) );
  XOR2_X1 U471 ( .A(G29GAT), .B(G43GAT), .Z(n405) );
  XNOR2_X1 U472 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n449) );
  XOR2_X1 U474 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n407) );
  XNOR2_X1 U475 ( .A(G106GAT), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n407), .B(n406), .ZN(n413) );
  XOR2_X1 U477 ( .A(KEYINPUT9), .B(n408), .Z(n411) );
  XNOR2_X1 U478 ( .A(G218GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n413), .B(n412), .ZN(n415) );
  AND2_X1 U481 ( .A1(G232GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n417) );
  INV_X1 U483 ( .A(KEYINPUT82), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n420) );
  XNOR2_X1 U485 ( .A(G99GAT), .B(G85GAT), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n418), .B(KEYINPUT71), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n432), .B(KEYINPUT80), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n449), .B(n421), .ZN(n424) );
  INV_X1 U490 ( .A(n422), .ZN(n423) );
  XOR2_X1 U491 ( .A(n424), .B(n423), .Z(n566) );
  XNOR2_X1 U492 ( .A(KEYINPUT36), .B(KEYINPUT106), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n566), .B(n425), .ZN(n596) );
  NOR2_X1 U494 ( .A1(n426), .A2(n596), .ZN(n429) );
  AND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n442) );
  XOR2_X1 U497 ( .A(n436), .B(n435), .Z(n440) );
  XOR2_X1 U498 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n438) );
  XNOR2_X1 U499 ( .A(KEYINPUT72), .B(KEYINPUT76), .ZN(n437) );
  XOR2_X1 U500 ( .A(n438), .B(n437), .Z(n439) );
  XOR2_X1 U501 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n444) );
  XNOR2_X1 U502 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n587) );
  XOR2_X1 U506 ( .A(n449), .B(KEYINPUT30), .Z(n451) );
  NAND2_X1 U507 ( .A1(G229GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n467) );
  XOR2_X1 U509 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n453) );
  XNOR2_X1 U510 ( .A(G8GAT), .B(G1GAT), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n465) );
  XOR2_X1 U512 ( .A(G141GAT), .B(G22GAT), .Z(n455) );
  XNOR2_X1 U513 ( .A(G36GAT), .B(G50GAT), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n455), .B(n454), .ZN(n463) );
  XOR2_X1 U515 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n457) );
  XNOR2_X1 U516 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(n461) );
  XOR2_X1 U518 ( .A(G113GAT), .B(G15GAT), .Z(n459) );
  XNOR2_X1 U519 ( .A(G169GAT), .B(G197GAT), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U521 ( .A(n461), .B(n460), .Z(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U523 ( .A(n465), .B(n464), .Z(n466) );
  XOR2_X1 U524 ( .A(n467), .B(n466), .Z(n554) );
  NOR2_X1 U525 ( .A1(n587), .A2(n554), .ZN(n496) );
  NAND2_X1 U526 ( .A1(n524), .A2(n496), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT38), .ZN(n511) );
  NOR2_X1 U528 ( .A1(n511), .A2(n540), .ZN(n471) );
  INV_X1 U529 ( .A(n554), .ZN(n582) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT46), .ZN(n473) );
  INV_X1 U531 ( .A(n566), .ZN(n547) );
  NOR2_X1 U532 ( .A1(n473), .A2(n547), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n563), .A2(n474), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT47), .ZN(n482) );
  NOR2_X1 U535 ( .A1(n596), .A2(n563), .ZN(n477) );
  INV_X1 U536 ( .A(KEYINPUT45), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n480) );
  INV_X1 U538 ( .A(n587), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n554), .A2(n478), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n481) );
  NOR2_X1 U541 ( .A1(n482), .A2(n481), .ZN(n483) );
  NOR2_X1 U542 ( .A1(n527), .A2(n534), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT54), .ZN(n579) );
  INV_X1 U544 ( .A(n485), .ZN(n486) );
  AND2_X1 U545 ( .A1(n578), .A2(n486), .ZN(n487) );
  AND2_X1 U546 ( .A1(n579), .A2(n487), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT55), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n540), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT120), .B(n490), .ZN(n575) );
  NAND2_X1 U550 ( .A1(n575), .A2(n547), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n547), .A2(n563), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT16), .B(n493), .Z(n494) );
  NOR2_X1 U553 ( .A1(n495), .A2(n494), .ZN(n514) );
  NAND2_X1 U554 ( .A1(n496), .A2(n514), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT102), .B(n497), .ZN(n505) );
  NOR2_X1 U556 ( .A1(n578), .A2(n505), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT34), .B(n498), .Z(n499) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  XNOR2_X1 U559 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n501) );
  NOR2_X1 U560 ( .A1(n527), .A2(n505), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1325GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n540), .A2(n505), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n504), .ZN(G1326GAT) );
  NOR2_X1 U566 ( .A1(n538), .A2(n505), .ZN(n506) );
  XOR2_X1 U567 ( .A(G22GAT), .B(n506), .Z(G1327GAT) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT39), .ZN(n509) );
  NOR2_X1 U570 ( .A1(n578), .A2(n511), .ZN(n508) );
  XOR2_X1 U571 ( .A(n509), .B(n508), .Z(G1328GAT) );
  NOR2_X1 U572 ( .A1(n527), .A2(n511), .ZN(n510) );
  XOR2_X1 U573 ( .A(G36GAT), .B(n510), .Z(G1329GAT) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n513) );
  NOR2_X1 U575 ( .A1(n538), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1331GAT) );
  INV_X1 U577 ( .A(n572), .ZN(n558) );
  NOR2_X1 U578 ( .A1(n582), .A2(n558), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n525), .A2(n514), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n578), .A2(n520), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(G57GAT), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U584 ( .A1(n527), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n518), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n540), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n538), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U591 ( .A(G78GAT), .B(n523), .Z(G1335GAT) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U593 ( .A1(n578), .A2(n531), .ZN(n526) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n526), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n531), .ZN(n528) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n540), .A2(n531), .ZN(n529) );
  XOR2_X1 U598 ( .A(KEYINPUT112), .B(n529), .Z(n530) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  NOR2_X1 U600 ( .A1(n538), .A2(n531), .ZN(n532) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n532), .Z(n533) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(KEYINPUT113), .B(n537), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n538), .A2(n553), .ZN(n539) );
  NOR2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n582), .A2(n548), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n543) );
  NAND2_X1 U610 ( .A1(n548), .A2(n572), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n592), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT115), .Z(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n553), .A2(n577), .ZN(n565) );
  NOR2_X1 U622 ( .A1(n554), .A2(n565), .ZN(n555) );
  XOR2_X1 U623 ( .A(G141GAT), .B(n555), .Z(G1344GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n558), .A2(n565), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U630 ( .A(n562), .B(n561), .Z(G1345GAT) );
  NOR2_X1 U631 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n582), .A2(n575), .ZN(n568) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(n568), .ZN(G1348GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n569) );
  XNOR2_X1 U639 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U640 ( .A(KEYINPUT56), .B(n571), .Z(n574) );
  NAND2_X1 U641 ( .A1(n572), .A2(n575), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NAND2_X1 U643 ( .A1(n575), .A2(n592), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT123), .Z(n584) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n594) );
  NAND2_X1 U648 ( .A1(n594), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n589) );
  NAND2_X1 U653 ( .A1(n594), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n591) );
  XOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT124), .Z(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NAND2_X1 U657 ( .A1(n594), .A2(n592), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n593), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U659 ( .A(n594), .ZN(n595) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U661 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(n599) );
  XOR2_X1 U663 ( .A(G218GAT), .B(n599), .Z(G1355GAT) );
endmodule

