//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n210), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n218), .B1(KEYINPUT1), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT68), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT69), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT70), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n214), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n206), .A2(G33), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT72), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT11), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT12), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G68), .ZN(new_n260));
  INV_X1    g0060(.A(new_n259), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(KEYINPUT12), .A3(new_n254), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n249), .B1(G1), .B2(new_n206), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n262), .C1(new_n263), .C2(new_n254), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n256), .B2(KEYINPUT11), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT14), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT13), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AND2_X1   g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n205), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n272), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G238), .A3(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G232), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n284), .B1(G226), .B2(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G97), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n279), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n269), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n279), .B1(new_n287), .B2(new_n288), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n281), .A2(new_n293), .A3(KEYINPUT13), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n268), .B(G169), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n282), .A2(new_n291), .A3(new_n269), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT13), .B1(new_n281), .B2(new_n293), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n297), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n268), .B1(new_n300), .B2(G169), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT75), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(G169), .B1(new_n292), .B2(new_n294), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT14), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT75), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n298), .A4(new_n295), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n267), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n296), .B2(new_n297), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n310), .A2(new_n266), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT78), .ZN(new_n316));
  INV_X1    g0116(.A(G226), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G1698), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(G223), .B2(G1698), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n285), .A2(new_n286), .ZN(new_n320));
  INV_X1    g0120(.A(G33), .ZN(new_n321));
  INV_X1    g0121(.A(G87), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n319), .A2(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n279), .A2(new_n274), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(new_n290), .B1(new_n324), .B2(G232), .ZN(new_n325));
  AOI21_X1  g0125(.A(G200), .B1(new_n325), .B2(new_n278), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n279), .A2(G232), .A3(new_n274), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n321), .A2(new_n322), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G223), .A2(G1698), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n317), .B2(G1698), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n321), .ZN(new_n332));
  NAND2_X1  g0132(.A1(KEYINPUT3), .A2(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n328), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n278), .B(new_n327), .C1(new_n335), .C2(new_n279), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(G190), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n316), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n311), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n323), .A2(new_n290), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n340), .A2(new_n309), .A3(new_n278), .A4(new_n327), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(KEYINPUT78), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  XOR2_X1   g0144(.A(KEYINPUT8), .B(G58), .Z(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n249), .C1(G1), .C2(new_n206), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT8), .B(G58), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n261), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(KEYINPUT77), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT77), .B1(new_n346), .B2(new_n348), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT16), .ZN(new_n353));
  INV_X1    g0153(.A(G58), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n254), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G58), .A2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n253), .A2(G159), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n332), .A2(new_n206), .A3(new_n333), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n333), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n254), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT76), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n360), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI211_X1 g0167(.A(KEYINPUT76), .B(new_n254), .C1(new_n363), .C2(new_n364), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n353), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n365), .A2(new_n359), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n249), .B1(new_n370), .B2(KEYINPUT16), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n352), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n343), .A2(new_n344), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n344), .B1(new_n343), .B2(new_n372), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n336), .A2(G169), .ZN(new_n376));
  INV_X1    g0176(.A(G179), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n336), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT18), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n352), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n320), .B2(new_n206), .ZN(new_n382));
  INV_X1    g0182(.A(new_n364), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n359), .B1(new_n384), .B2(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n365), .A2(new_n366), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n248), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n381), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n378), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n375), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G50), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n261), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G150), .ZN(new_n398));
  INV_X1    g0198(.A(new_n253), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n398), .A2(new_n399), .B1(new_n201), .B2(new_n206), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n251), .B2(new_n345), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n397), .B1(new_n396), .B2(new_n263), .C1(new_n401), .C2(new_n249), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT9), .ZN(new_n403));
  INV_X1    g0203(.A(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G222), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n334), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n290), .C1(G77), .C2(new_n334), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n324), .A2(G226), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n278), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G200), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n309), .B2(new_n410), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n403), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(KEYINPUT74), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT10), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n403), .A2(new_n416), .A3(new_n413), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n410), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n402), .B(new_n422), .C1(G179), .C2(new_n410), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT15), .B(G87), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n250), .B1(new_n206), .B2(new_n202), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n347), .A2(new_n399), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n248), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g0228(.A(new_n428), .B(KEYINPUT73), .Z(new_n429));
  MUX2_X1   g0229(.A(new_n259), .B(new_n263), .S(G77), .Z(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G238), .A2(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n334), .B(new_n433), .C1(new_n283), .C2(G1698), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n290), .C1(G107), .C2(new_n334), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n324), .A2(G244), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n278), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n421), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(G179), .B2(new_n437), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(G200), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n309), .B2(new_n437), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OR4_X1    g0245(.A1(new_n315), .A2(new_n395), .A3(new_n424), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n404), .A2(G257), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G264), .A2(G1698), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n334), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G303), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n320), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n290), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  INV_X1    g0258(.A(G41), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G270), .A3(new_n279), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT86), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT86), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n461), .A2(new_n464), .A3(G270), .A4(new_n279), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n273), .A2(new_n456), .A3(new_n458), .A4(new_n460), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT87), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n461), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n462), .A2(KEYINPUT86), .B1(new_n470), .B2(new_n273), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT87), .B1(new_n471), .B2(new_n465), .ZN(new_n472));
  OAI211_X1 g0272(.A(G190), .B(new_n453), .C1(new_n469), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  INV_X1    g0274(.A(G97), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n474), .B(new_n206), .C1(G33), .C2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n248), .C1(new_n206), .C2(G116), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT20), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n261), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n249), .B(new_n259), .C1(G1), .C2(new_n321), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n479), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n453), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n467), .A2(new_n468), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(KEYINPUT87), .A3(new_n465), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n473), .B(new_n483), .C1(new_n311), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  OAI21_X1  g0289(.A(G169), .B1(new_n478), .B2(new_n482), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n483), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(G179), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n453), .B1(new_n469), .B2(new_n472), .ZN(new_n494));
  INV_X1    g0294(.A(new_n490), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(KEYINPUT21), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n488), .A2(new_n491), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(G1698), .B1(new_n332), .B2(new_n333), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT90), .A3(G250), .ZN(new_n499));
  OAI211_X1 g0299(.A(G250), .B(new_n404), .C1(new_n285), .C2(new_n286), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT90), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G257), .A2(G1698), .ZN(new_n504));
  INV_X1    g0304(.A(G294), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n320), .A2(new_n504), .B1(new_n321), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n290), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n461), .A2(G264), .A3(new_n279), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n507), .A2(new_n377), .A3(new_n466), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n499), .B2(new_n502), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n466), .B(new_n508), .C1(new_n510), .C2(new_n279), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n421), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n206), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n334), .A2(new_n515), .A3(new_n206), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OR3_X1    g0317(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT88), .B1(new_n519), .B2(G20), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n519), .A2(KEYINPUT88), .A3(G20), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT24), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n517), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n249), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n481), .ZN(new_n530));
  INV_X1    g0330(.A(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n261), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  AOI22_X1  g0336(.A1(G107), .A2(new_n530), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n509), .B(new_n512), .C1(new_n529), .C2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n507), .A2(G190), .A3(new_n466), .A4(new_n508), .ZN(new_n540));
  INV_X1    g0340(.A(new_n528), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n527), .B1(new_n517), .B2(new_n524), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n248), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n511), .A2(G200), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n540), .A2(new_n543), .A3(new_n544), .A4(new_n537), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n261), .A2(new_n475), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n481), .B2(new_n475), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT6), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n550), .A2(new_n475), .A3(G107), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n531), .B1(new_n363), .B2(new_n364), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n548), .B1(new_n558), .B2(new_n248), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n461), .A2(G257), .A3(new_n279), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n466), .ZN(new_n561));
  OAI211_X1 g0361(.A(G244), .B(new_n404), .C1(new_n285), .C2(new_n286), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT79), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n563), .A2(KEYINPUT4), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n474), .ZN(new_n567));
  INV_X1    g0367(.A(G250), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n404), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n334), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n334), .A2(G244), .A3(new_n404), .A4(new_n564), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n561), .B1(new_n290), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n573), .B2(KEYINPUT81), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n290), .ZN(new_n576));
  INV_X1    g0376(.A(new_n561), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n576), .A2(KEYINPUT81), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n559), .B(new_n574), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n377), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT82), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n577), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n421), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n573), .A2(new_n584), .A3(new_n377), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n552), .B1(new_n550), .B2(new_n549), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n586), .A2(new_n206), .B1(new_n202), .B2(new_n399), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n248), .B1(new_n587), .B2(new_n556), .ZN(new_n588));
  INV_X1    g0388(.A(new_n548), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n581), .A2(new_n583), .A3(new_n585), .A4(new_n590), .ZN(new_n591));
  XOR2_X1   g0391(.A(KEYINPUT15), .B(G87), .Z(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n259), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n322), .A2(new_n475), .A3(new_n531), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n288), .A2(new_n206), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT19), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n206), .B(G68), .C1(new_n285), .C2(new_n286), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n250), .B2(new_n475), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(KEYINPUT85), .B(new_n593), .C1(new_n248), .C2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT85), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n248), .ZN(new_n603));
  INV_X1    g0403(.A(new_n593), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n601), .A2(new_n605), .B1(new_n425), .B2(new_n481), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n334), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n498), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n279), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OR3_X1    g0413(.A1(new_n458), .A2(KEYINPUT83), .A3(new_n568), .ZN(new_n614));
  AND2_X1   g0414(.A1(KEYINPUT83), .A2(G250), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n458), .B1(new_n615), .B2(G274), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n290), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n421), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n334), .A2(G238), .A3(new_n404), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n519), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n609), .B2(new_n610), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n377), .B(new_n619), .C1(new_n622), .C2(new_n279), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n606), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n593), .B1(new_n600), .B2(new_n248), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(new_n602), .ZN(new_n626));
  OAI211_X1 g0426(.A(G190), .B(new_n619), .C1(new_n622), .C2(new_n279), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n530), .A2(G87), .ZN(new_n628));
  OAI21_X1  g0428(.A(G200), .B1(new_n613), .B2(new_n617), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n579), .A2(new_n591), .A3(new_n624), .A4(new_n630), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n497), .A2(new_n546), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n447), .A2(new_n632), .ZN(G372));
  NAND2_X1  g0433(.A1(new_n314), .A2(new_n440), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n375), .B1(new_n308), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT92), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n391), .B1(new_n390), .B2(new_n378), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n372), .A2(KEYINPUT18), .A3(new_n379), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n380), .A2(new_n392), .A3(KEYINPUT92), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n420), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n496), .A2(new_n491), .A3(new_n493), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT91), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n496), .A2(new_n491), .A3(KEYINPUT91), .A4(new_n493), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n539), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n631), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n545), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n624), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n624), .A2(new_n630), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n591), .ZN(new_n654));
  INV_X1    g0454(.A(new_n591), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(KEYINPUT26), .A3(new_n624), .A4(new_n630), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n423), .B(new_n642), .C1(new_n446), .C2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(new_n539), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT93), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n529), .B2(new_n538), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n539), .A2(new_n545), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT94), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(KEYINPUT94), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n666), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n643), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n675), .A2(new_n678), .B1(new_n660), .B2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n645), .A2(new_n646), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n483), .A2(new_n676), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n497), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n209), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n594), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n216), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n658), .A2(KEYINPUT29), .A3(new_n666), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n483), .B1(new_n487), .B2(new_n311), .ZN(new_n697));
  INV_X1    g0497(.A(new_n473), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n643), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n631), .A2(new_n546), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n676), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT31), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n613), .A2(new_n617), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n704), .A2(G179), .A3(new_n573), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n494), .A3(new_n511), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n704), .A2(new_n508), .A3(new_n507), .A4(new_n573), .ZN(new_n707));
  OAI211_X1 g0507(.A(G179), .B(new_n453), .C1(new_n469), .C2(new_n472), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n487), .A2(new_n710), .A3(G179), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n707), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n706), .B1(new_n712), .B2(KEYINPUT30), .ZN(new_n713));
  INV_X1    g0513(.A(new_n707), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n710), .B1(new_n487), .B2(G179), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n666), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n703), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n666), .C1(new_n713), .C2(new_n719), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n696), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n648), .B(new_n545), .C1(new_n660), .C2(new_n643), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n657), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n676), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n695), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n694), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n690), .A2(G1), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n685), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n683), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n683), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n214), .B1(G20), .B2(new_n421), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n206), .A2(new_n377), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G190), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n206), .A2(G179), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n309), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n746), .A2(new_n747), .B1(new_n750), .B2(G283), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G20), .A3(new_n309), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n334), .B1(new_n754), .B2(G329), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n751), .B(new_n755), .C1(new_n451), .C2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n744), .B(KEYINPUT98), .Z(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n745), .A2(new_n309), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G326), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n761), .A2(new_n762), .B1(new_n505), .B2(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n759), .A2(G311), .B1(new_n766), .B2(KEYINPUT100), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(KEYINPUT100), .B2(new_n766), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT101), .Z(new_n769));
  NOR3_X1   g0569(.A1(new_n758), .A2(new_n309), .A3(G200), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n757), .B(new_n769), .C1(G322), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n756), .A2(new_n322), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(G107), .B2(new_n750), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G50), .A2(new_n760), .B1(new_n746), .B2(G68), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n753), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n773), .B(new_n774), .C1(new_n777), .C2(KEYINPUT99), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n320), .B1(new_n764), .B2(G97), .ZN(new_n779));
  INV_X1    g0579(.A(new_n770), .ZN(new_n780));
  INV_X1    g0580(.A(new_n759), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n779), .B1(new_n780), .B2(new_n354), .C1(new_n202), .C2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n778), .B(new_n782), .C1(KEYINPUT99), .C2(new_n777), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n743), .B1(new_n771), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n740), .A2(new_n743), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n688), .A2(new_n334), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n241), .A2(new_n457), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT96), .Z(new_n790));
  AOI211_X1 g0590(.A(new_n788), .B(new_n790), .C1(new_n457), .C2(new_n217), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n209), .A2(new_n334), .ZN(new_n792));
  INV_X1    g0592(.A(G355), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n792), .A2(new_n793), .B1(G116), .B2(new_n209), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n786), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n742), .A2(new_n784), .A3(new_n735), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n737), .A2(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n440), .A2(new_n676), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n443), .B1(new_n431), .B2(new_n666), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n440), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n658), .B2(new_n666), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n444), .A2(new_n676), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n650), .B2(new_n657), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n735), .B1(new_n805), .B2(new_n724), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n724), .B2(new_n805), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G137), .A2(new_n760), .B1(new_n746), .B2(G150), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n780), .B2(new_n809), .C1(new_n775), .C2(new_n781), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  AOI21_X1  g0611(.A(new_n320), .B1(new_n754), .B2(G132), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n254), .B2(new_n749), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n765), .A2(new_n354), .B1(new_n756), .B2(new_n396), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n760), .A2(G303), .B1(new_n750), .B2(G87), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n531), .B2(new_n756), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n320), .B1(new_n818), .B2(new_n753), .C1(new_n765), .C2(new_n475), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n759), .B2(G116), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n505), .B2(new_n780), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n746), .A2(KEYINPUT102), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n746), .A2(KEYINPUT102), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n817), .B(new_n821), .C1(G283), .C2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n743), .B1(new_n815), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n743), .A2(new_n738), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n734), .B1(new_n202), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n800), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n739), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n807), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n732), .A2(new_n205), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT106), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n267), .A2(new_n676), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n307), .A2(new_n313), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n836), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n302), .B2(new_n306), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n830), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n721), .B2(new_n722), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n343), .A2(new_n372), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n370), .A2(KEYINPUT16), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n389), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n346), .A2(new_n348), .ZN(new_n846));
  INV_X1    g0646(.A(new_n664), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n845), .A2(new_n846), .B1(new_n378), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n390), .A2(new_n378), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n390), .A2(new_n847), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n843), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n845), .A2(new_n846), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n847), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n637), .A2(new_n638), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n339), .A2(KEYINPUT78), .A3(new_n341), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT78), .B1(new_n339), .B2(new_n341), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT17), .B1(new_n862), .B2(new_n390), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n343), .A2(new_n344), .A3(new_n372), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n858), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n842), .B1(new_n856), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT38), .B(new_n855), .C1(new_n394), .C2(new_n858), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n835), .B(KEYINPUT40), .C1(new_n841), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT31), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n632), .B2(new_n676), .ZN(new_n872));
  INV_X1    g0672(.A(new_n706), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n717), .B2(new_n718), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n712), .A2(KEYINPUT30), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n676), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n722), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n308), .A2(new_n314), .A3(new_n838), .ZN(new_n878));
  INV_X1    g0678(.A(new_n839), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n800), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n869), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT106), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n870), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n373), .B2(new_n374), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n863), .A2(KEYINPUT104), .A3(new_n864), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(new_n639), .A3(new_n640), .A4(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n852), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT105), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n843), .A2(new_n851), .A3(new_n852), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n854), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT105), .B1(new_n888), .B2(new_n889), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n842), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n868), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n717), .A2(new_n718), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n875), .A3(new_n706), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n666), .A2(new_n899), .B1(new_n702), .B2(KEYINPUT31), .ZN(new_n900));
  INV_X1    g0700(.A(new_n722), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n882), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n884), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n447), .A2(new_n877), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT107), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n696), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  INV_X1    g0708(.A(new_n868), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n308), .A2(new_n666), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n867), .A2(new_n868), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n837), .A2(new_n839), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n798), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n803), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n920), .B2(KEYINPUT103), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(KEYINPUT103), .B2(new_n920), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n641), .A2(new_n664), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n915), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n446), .B1(new_n695), .B2(new_n728), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n642), .A2(new_n423), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n924), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n834), .B1(new_n908), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n908), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(G116), .A3(new_n215), .A4(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n355), .A2(new_n216), .A3(new_n202), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n254), .A2(G50), .ZN(new_n936));
  OAI211_X1 g0736(.A(G1), .B(new_n731), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  NAND2_X1  g0738(.A1(new_n655), .A2(new_n666), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT108), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n579), .B(new_n591), .C1(new_n559), .C2(new_n676), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n660), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n666), .B1(new_n943), .B2(new_n591), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n675), .A2(new_n678), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n942), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n947), .B2(KEYINPUT42), .ZN(new_n948));
  INV_X1    g0748(.A(new_n942), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n945), .A2(KEYINPUT42), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n626), .A2(new_n628), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n651), .A2(new_n952), .A3(new_n666), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n666), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n624), .A3(new_n630), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n686), .A2(new_n949), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n948), .A2(new_n958), .A3(new_n957), .A4(new_n950), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n961), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n689), .B(KEYINPUT41), .Z(new_n967));
  NAND3_X1  g0767(.A1(new_n673), .A2(new_n674), .A3(new_n677), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n684), .B1(new_n946), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n945), .A2(new_n685), .A3(new_n968), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n729), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n686), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n660), .A2(new_n676), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n945), .A2(new_n976), .A3(new_n942), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n945), .A2(new_n976), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT44), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n949), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT44), .B1(new_n679), .B2(new_n942), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n975), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n979), .A2(new_n980), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n686), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n974), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n967), .B1(new_n991), .B2(new_n729), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n733), .A2(G1), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n966), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n785), .B1(new_n209), .B2(new_n425), .C1(new_n231), .C2(new_n788), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n995), .A2(new_n735), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n320), .B1(new_n753), .B2(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n761), .A2(new_n818), .B1(new_n749), .B2(new_n475), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G107), .C2(new_n764), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G283), .A2(new_n759), .B1(new_n770), .B2(G303), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n756), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(G116), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT46), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n825), .A2(G294), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1001), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G50), .A2(new_n759), .B1(new_n770), .B2(G150), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1002), .A2(G58), .B1(new_n754), .B2(G137), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n760), .A2(G143), .B1(G68), .B2(new_n764), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n334), .B1(new_n749), .B2(new_n202), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT109), .Z(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n775), .B2(new_n824), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1006), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT47), .Z(new_n1015));
  INV_X1    g0815(.A(new_n743), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n996), .B1(new_n741), .B2(new_n956), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n994), .A2(new_n1017), .ZN(G387));
  NAND3_X1  g0818(.A1(new_n970), .A2(new_n993), .A3(new_n971), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT110), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n688), .A2(new_n531), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n457), .B1(new_n254), .B2(new_n202), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n691), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n347), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n787), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n236), .A2(new_n457), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1021), .B1(new_n691), .B2(new_n792), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n734), .B1(new_n1030), .B2(new_n786), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n764), .A2(new_n592), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n780), .B2(new_n396), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT113), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n760), .A2(G159), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT112), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n334), .B1(new_n753), .B2(new_n398), .C1(new_n749), .C2(new_n475), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n746), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1038), .A2(new_n347), .B1(new_n202), .B2(new_n756), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(new_n759), .C2(G68), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1034), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n320), .B1(new_n753), .B2(new_n762), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n770), .A2(G317), .B1(G322), .B2(new_n760), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n451), .B2(new_n781), .C1(new_n818), .C2(new_n824), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1002), .A2(G294), .B1(new_n764), .B2(G283), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1042), .B(new_n1051), .C1(G116), .C2(new_n750), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1041), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1031), .B1(new_n675), .B2(new_n741), .C1(new_n1054), .C2(new_n1016), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1020), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n974), .A2(new_n690), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n729), .B2(new_n972), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(G393));
  NAND3_X1  g0859(.A1(new_n987), .A2(new_n993), .A3(new_n990), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n787), .A2(new_n244), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n740), .B(new_n743), .C1(new_n688), .C2(G97), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n734), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n334), .B1(new_n754), .B2(G322), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n531), .B2(new_n749), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n770), .A2(G311), .B1(G317), .B2(new_n760), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(G283), .C2(new_n1002), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n759), .A2(G294), .B1(G116), .B2(new_n764), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n451), .B2(new_n824), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT115), .Z(new_n1071));
  OAI221_X1 g0871(.A(new_n334), .B1(new_n749), .B2(new_n322), .C1(new_n765), .C2(new_n202), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n756), .A2(new_n254), .B1(new_n809), .B2(new_n753), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n825), .A2(G50), .B1(KEYINPUT114), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT114), .B2(new_n1073), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1072), .B(new_n1075), .C1(new_n345), .C2(new_n759), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n770), .A2(G159), .B1(G150), .B2(new_n760), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  AOI22_X1  g0878(.A1(new_n1068), .A2(new_n1071), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1063), .B1(new_n942), .B2(new_n741), .C1(new_n1016), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1060), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n981), .A2(new_n975), .A3(new_n986), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n686), .B1(new_n988), .B2(new_n989), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n690), .B1(new_n1084), .B2(new_n974), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n973), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(G390));
  NAND2_X1  g0888(.A1(new_n723), .A2(new_n880), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n914), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n920), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n911), .A2(new_n912), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n443), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n431), .A2(new_n666), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n440), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n798), .B1(new_n727), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n914), .B1(new_n1097), .B2(new_n918), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n897), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1093), .A2(KEYINPUT116), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT116), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1090), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1089), .B1(new_n1103), .B2(KEYINPUT116), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n918), .B1(new_n723), .B2(new_n830), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1090), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1097), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n803), .A2(new_n919), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n724), .A2(new_n446), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n925), .A2(new_n926), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT117), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n690), .B1(new_n1105), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT117), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n911), .A2(new_n738), .A3(new_n912), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n345), .A2(new_n743), .A3(new_n738), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n770), .A2(G116), .B1(G77), .B2(new_n764), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT119), .Z(new_n1124));
  AOI211_X1 g0924(.A(new_n334), .B(new_n772), .C1(G294), .C2(new_n754), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n760), .A2(G283), .B1(new_n750), .B2(G68), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n475), .B2(new_n781), .C1(new_n531), .C2(new_n824), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT54), .B(G143), .Z(new_n1129));
  AOI22_X1  g0929(.A1(G132), .A2(new_n770), .B1(new_n759), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n334), .B1(new_n753), .B2(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n765), .A2(new_n775), .B1(new_n749), .B2(new_n396), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G128), .C2(new_n760), .ZN(new_n1134));
  INV_X1    g0934(.A(G137), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1130), .B(new_n1134), .C1(new_n1135), .C2(new_n824), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n756), .A2(new_n398), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT118), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1124), .A2(new_n1128), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n734), .B(new_n1122), .C1(new_n1140), .C2(new_n743), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n993), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(new_n1105), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1120), .A2(new_n1145), .ZN(G378));
  NAND3_X1  g0946(.A1(new_n1102), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1113), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n424), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1149), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n420), .A2(new_n423), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n402), .A2(new_n847), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1150), .A2(new_n402), .A3(new_n847), .A4(new_n1152), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n888), .A2(new_n889), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT105), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n893), .A3(new_n890), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n909), .B1(new_n1162), .B2(new_n842), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n841), .A2(KEYINPUT40), .ZN(new_n1164));
  OAI21_X1  g0964(.A(G330), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1158), .B1(new_n884), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n915), .A2(new_n922), .A3(new_n923), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n882), .B1(new_n902), .B2(new_n916), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n835), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n881), .A2(KEYINPUT106), .A3(new_n882), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1155), .A2(KEYINPUT122), .A3(new_n1156), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT122), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n696), .B1(new_n897), .B2(new_n903), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1171), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1166), .A2(new_n1167), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1167), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1148), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1148), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n689), .A3(new_n1183), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n884), .A2(new_n1165), .A3(new_n1174), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1157), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n924), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1166), .A2(new_n1167), .A3(new_n1177), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n993), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n734), .B1(new_n396), .B2(new_n828), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT121), .ZN(new_n1191));
  INV_X1    g0991(.A(G283), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n765), .A2(new_n254), .B1(new_n1192), .B2(new_n753), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n781), .A2(new_n425), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G107), .C2(new_n770), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n760), .A2(G116), .B1(new_n750), .B2(G58), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n475), .B2(new_n1038), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT120), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n459), .B(new_n320), .C1(new_n756), .C2(new_n202), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1195), .B(new_n1200), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT58), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n396), .B1(new_n285), .B2(G41), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G128), .A2(new_n770), .B1(new_n759), .B2(G137), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G125), .A2(new_n760), .B1(new_n746), .B2(G132), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1002), .A2(new_n1129), .B1(new_n764), .B2(G150), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n750), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1202), .B(new_n1203), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1191), .B1(new_n1214), .B2(new_n743), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1175), .B2(new_n739), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1189), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1184), .A2(new_n1217), .ZN(G375));
  INV_X1    g1018(.A(new_n1111), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1113), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n967), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1116), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n734), .B1(new_n254), .B2(new_n828), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n320), .B1(new_n754), .B2(G128), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n354), .B2(new_n749), .C1(new_n780), .C2(new_n1135), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G150), .B2(new_n759), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n760), .A2(G132), .B1(G50), .B2(new_n764), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n775), .B2(new_n756), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n825), .B2(new_n1129), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n531), .A2(new_n781), .B1(new_n780), .B2(new_n1192), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1032), .B1(new_n451), .B2(new_n753), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n761), .A2(new_n505), .B1(new_n475), .B2(new_n756), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT123), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n334), .B1(new_n750), .B2(G77), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n824), .A2(new_n479), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1227), .A2(new_n1230), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1224), .B1(new_n1239), .B2(new_n1016), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n917), .B2(new_n738), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1111), .B2(new_n993), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1223), .A2(new_n1242), .ZN(G381));
  XNOR2_X1  g1043(.A(G375), .B(KEYINPUT124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n994), .A2(new_n1087), .A3(new_n1017), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1056), .A2(new_n1058), .A3(new_n796), .A4(new_n737), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G384), .A2(new_n1245), .A3(G381), .A4(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1244), .A2(new_n1247), .A3(G378), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n665), .A2(G213), .ZN(new_n1249));
  OR3_X1    g1049(.A1(new_n1244), .A2(G378), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(G407), .A2(new_n1250), .A3(G213), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1189), .A2(new_n1216), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1113), .B2(new_n1147), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1255), .B2(new_n1222), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1252), .B1(new_n1256), .B2(G378), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1183), .A2(new_n689), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1217), .C1(new_n1258), .C2(new_n1181), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1148), .A2(new_n1180), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1217), .B1(new_n1260), .B2(new_n967), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1144), .B1(new_n1119), .B2(new_n1115), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(KEYINPUT125), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1257), .A2(new_n1259), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n689), .B(new_n1116), .C1(new_n1221), .C2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT60), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1242), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n832), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G384), .B(new_n1242), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1264), .A2(new_n1249), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT126), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1264), .A2(new_n1249), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n665), .A2(G213), .A3(G2897), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1269), .A2(new_n1270), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1264), .A2(new_n1249), .A3(new_n1272), .A4(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1276), .A2(new_n1282), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1287), .A2(new_n1246), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n994), .A2(new_n1087), .A3(new_n1017), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1087), .B1(new_n994), .B2(new_n1017), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G387), .A2(G390), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1287), .A2(new_n1246), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1245), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1286), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1297), .B2(new_n1273), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1264), .A2(KEYINPUT63), .A3(new_n1249), .A4(new_n1272), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1283), .A3(new_n1299), .A4(new_n1282), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1262), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1271), .A3(new_n1259), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G378), .B1(new_n1184), .B2(new_n1217), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1259), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1272), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1303), .A2(new_n1295), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1295), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  AOI211_X1 g1110(.A(KEYINPUT127), .B(new_n1295), .C1(new_n1306), .C2(new_n1303), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


