//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n591, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n460));
  XOR2_X1   g035(.A(KEYINPUT67), .B(G2105), .Z(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n463), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n462), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n459), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n459), .A2(new_n463), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n477), .A2(G124), .B1(new_n479), .B2(G136), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n485));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n471), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n461), .A2(new_n490), .A3(G138), .A4(new_n459), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(G164));
  AND2_X1   g067(.A1(KEYINPUT6), .A2(G651), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT6), .A2(G651), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G50), .ZN(new_n497));
  INV_X1    g072(.A(G88), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n499), .A2(new_n500), .B1(new_n493), .B2(new_n494), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT68), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n502), .A2(new_n510), .ZN(G166));
  NOR2_X1   g086(.A1(new_n493), .A2(new_n494), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G51), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n495), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n500), .A2(new_n499), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n515), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G168));
  INV_X1    g099(.A(new_n501), .ZN(new_n525));
  AOI22_X1  g100(.A1(G90), .A2(new_n525), .B1(new_n514), .B2(G52), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n503), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(G171));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G56), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n519), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n503), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(new_n535), .B2(new_n534), .ZN(new_n537));
  AOI22_X1  g112(.A1(G81), .A2(new_n525), .B1(new_n514), .B2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n514), .A2(G53), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(KEYINPUT72), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n546), .B(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n503), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n525), .A2(G91), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(G299));
  NAND2_X1  g128(.A1(new_n528), .A2(new_n530), .ZN(G301));
  AND2_X1   g129(.A1(new_n522), .A2(new_n523), .ZN(G286));
  INV_X1    g130(.A(G166), .ZN(G303));
  INV_X1    g131(.A(G74), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n503), .B1(new_n519), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(G49), .B2(new_n514), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n525), .A2(G87), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(G288));
  OAI211_X1 g136(.A(G48), .B(G543), .C1(new_n493), .C2(new_n494), .ZN(new_n562));
  INV_X1    g137(.A(G86), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n501), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(G61), .B1(new_n500), .B2(new_n499), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n503), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G305));
  INV_X1    g144(.A(G47), .ZN(new_n570));
  INV_X1    g145(.A(G85), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n496), .A2(new_n570), .B1(new_n571), .B2(new_n501), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n503), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(new_n525), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT10), .Z(new_n578));
  NAND2_X1  g153(.A1(G79), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G66), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n519), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n514), .B2(G54), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(G171), .B2(new_n584), .ZN(G284));
  OAI21_X1  g161(.A(new_n585), .B1(G171), .B2(new_n584), .ZN(G321));
  NOR2_X1   g162(.A1(G299), .A2(G868), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g164(.A(new_n588), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g165(.A(new_n583), .ZN(new_n591));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n459), .A2(new_n464), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT12), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(G2100), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(G2100), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n477), .A2(G123), .ZN(new_n604));
  OAI221_X1 g179(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n461), .C2(G111), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n479), .A2(G135), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(G2096), .Z(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n603), .A3(new_n608), .ZN(G156));
  XOR2_X1   g184(.A(G1341), .B(G1348), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT74), .ZN(new_n611));
  XOR2_X1   g186(.A(G2451), .B(G2454), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT16), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n611), .B(new_n613), .Z(new_n614));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n615));
  XNOR2_X1  g190(.A(G2427), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(new_n617), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n614), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(G14), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT75), .Z(G401));
  XNOR2_X1  g201(.A(G2067), .B(G2678), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT76), .ZN(new_n628));
  NOR2_X1   g203(.A1(G2072), .A2(G2078), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n442), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2084), .B(G2090), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n628), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n628), .A2(new_n630), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n630), .B(KEYINPUT17), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n635), .B(new_n632), .C1(new_n628), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n628), .A3(new_n631), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2096), .B(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT77), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(G227));
  XOR2_X1   g217(.A(KEYINPUT78), .B(KEYINPUT19), .Z(new_n643));
  XNOR2_X1  g218(.A(G1971), .B(G1976), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1956), .B(G2474), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1961), .B(G1966), .Z(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT79), .Z(new_n651));
  AND2_X1   g226(.A1(new_n647), .A2(new_n648), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n645), .A2(new_n652), .A3(new_n649), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1991), .B(G1996), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G229));
  MUX2_X1   g237(.A(G23), .B(G288), .S(G16), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT33), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G22), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(G166), .B2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(G1971), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(G6), .A2(G16), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n568), .B2(G16), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT32), .B(G1981), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n667), .A2(new_n668), .A3(new_n673), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT82), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n669), .A2(G24), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT80), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G290), .B2(G16), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n477), .A2(G119), .B1(new_n479), .B2(G131), .ZN(new_n688));
  OAI221_X1 g263(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n461), .C2(G107), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(G25), .B(new_n690), .S(G29), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT35), .B(G1991), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  AOI211_X1 g269(.A(new_n687), .B(new_n694), .C1(KEYINPUT83), .C2(KEYINPUT36), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n681), .A2(new_n682), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G21), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G168), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT94), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT95), .B(G1966), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT96), .Z(new_n704));
  NOR2_X1   g279(.A1(G171), .A2(new_n669), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G5), .B2(new_n669), .ZN(new_n706));
  INV_X1    g281(.A(G1961), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT97), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT30), .B(G28), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OR2_X1    g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  NAND2_X1  g287(.A1(KEYINPUT31), .A2(G11), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n710), .A2(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n607), .B2(new_n711), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n701), .B2(new_n702), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n704), .A2(new_n709), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT98), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n696), .A2(new_n697), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n669), .A2(G20), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT23), .Z(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G299), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1956), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n711), .A2(G32), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n464), .A2(G105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT91), .ZN(new_n728));
  INV_X1    g303(.A(G141), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n478), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  INV_X1    g307(.A(G129), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n476), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n726), .B1(new_n735), .B2(new_n711), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g313(.A1(G160), .A2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n711), .B1(new_n740), .B2(G34), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(KEYINPUT89), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(G34), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n741), .B2(KEYINPUT89), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n739), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n736), .A2(new_n738), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n591), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G4), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n711), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n711), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT29), .Z(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n747), .B1(new_n749), .B2(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n725), .B(new_n755), .C1(new_n707), .C2(new_n706), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G19), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n540), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT84), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n753), .A2(new_n754), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT99), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n711), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n477), .A2(G128), .B1(new_n479), .B2(G140), .ZN(new_n765));
  NOR2_X1   g340(.A1(G104), .A2(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT85), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2067), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n749), .A2(new_n750), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  NAND2_X1  g349(.A1(G164), .A2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G27), .B2(G29), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n772), .B(new_n777), .C1(new_n774), .C2(new_n776), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n756), .A2(new_n760), .A3(new_n762), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n711), .A2(G33), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT25), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n479), .A2(G139), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n782), .B(new_n783), .C1(new_n461), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT86), .Z(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(new_n711), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G2072), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT87), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n745), .A2(new_n746), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n736), .A2(new_n738), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n787), .C2(G2072), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n789), .A2(KEYINPUT93), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT93), .B1(new_n789), .B2(new_n793), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n779), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n698), .A2(new_n719), .A3(new_n720), .A4(new_n796), .ZN(G150));
  INV_X1    g372(.A(G150), .ZN(G311));
  NAND2_X1  g373(.A1(new_n591), .A2(G559), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT38), .ZN(new_n800));
  AOI22_X1  g375(.A1(G93), .A2(new_n525), .B1(new_n514), .B2(G55), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n503), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n539), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n539), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n800), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n809), .A2(new_n810), .A3(G860), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n803), .A2(G860), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n813), .ZN(G145));
  NOR2_X1   g389(.A1(new_n786), .A2(new_n735), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n769), .B(G164), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n785), .B(KEYINPUT86), .ZN(new_n817));
  INV_X1    g392(.A(new_n735), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR3_X1    g394(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n477), .A2(G130), .B1(new_n479), .B2(G142), .ZN(new_n821));
  OAI221_X1 g396(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n599), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n690), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(KEYINPUT100), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n815), .B2(new_n819), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n825), .B(KEYINPUT100), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n820), .B2(new_n827), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n607), .B(G160), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n482), .ZN(new_n833));
  AOI21_X1  g408(.A(G37), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n833), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n828), .B2(new_n830), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT101), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(KEYINPUT101), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(G395));
  NAND2_X1  g416(.A1(new_n803), .A2(new_n584), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  NAND2_X1  g418(.A1(G299), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n549), .A2(KEYINPUT103), .A3(new_n551), .A4(new_n552), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n591), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n583), .A2(new_n843), .A3(G299), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n846), .A2(KEYINPUT41), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(new_n846), .B2(new_n847), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n807), .B(new_n594), .ZN(new_n853));
  MUX2_X1   g428(.A(new_n849), .B(new_n852), .S(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT42), .ZN(new_n855));
  XNOR2_X1  g430(.A(G166), .B(G288), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n575), .B(new_n568), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n855), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n842), .B1(new_n860), .B2(new_n584), .ZN(G295));
  OAI21_X1  g436(.A(new_n842), .B1(new_n860), .B2(new_n584), .ZN(G331));
  NOR2_X1   g437(.A1(G171), .A2(G168), .ZN(new_n863));
  NOR2_X1   g438(.A1(G286), .A2(G301), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n806), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(G286), .A2(G301), .ZN(new_n866));
  NAND2_X1  g441(.A1(G171), .A2(G168), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n807), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g445(.A(KEYINPUT104), .B(new_n806), .C1(new_n863), .C2(new_n864), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n848), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(new_n868), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n872), .A2(KEYINPUT105), .B1(new_n852), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n875), .A3(new_n859), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n874), .A2(new_n848), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n852), .A2(new_n870), .A3(new_n871), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n852), .A2(new_n870), .A3(KEYINPUT106), .A4(new_n871), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n859), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n876), .B(new_n877), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n876), .A2(new_n877), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n873), .A2(new_n875), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n858), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT43), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT44), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT43), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(G397));
  INV_X1    g473(.A(KEYINPUT54), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n489), .A2(new_n491), .ZN(new_n900));
  INV_X1    g475(.A(new_n487), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G1384), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(G164), .B2(G1384), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n473), .B(KEYINPUT123), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT53), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(G2078), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G40), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n908), .A2(new_n462), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G40), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n462), .A2(new_n913), .A3(new_n473), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n904), .A2(new_n906), .A3(new_n774), .A4(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n907), .A2(new_n912), .B1(new_n915), .B2(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n902), .A2(KEYINPUT109), .A3(new_n903), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(G164), .B2(G1384), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n902), .A2(new_n903), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n914), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n707), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n899), .B1(new_n926), .B2(G171), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT45), .B1(new_n917), .B2(new_n919), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n904), .A2(new_n914), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n930), .A2(new_n910), .B1(new_n909), .B2(new_n915), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(G301), .A3(new_n925), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n702), .B1(new_n928), .B2(new_n929), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n921), .A2(new_n746), .A3(new_n914), .A4(new_n923), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G8), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  NOR2_X1   g513(.A1(G168), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT51), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n934), .A2(KEYINPUT121), .A3(new_n935), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT121), .B1(new_n934), .B2(new_n935), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n942), .A2(new_n943), .A3(G286), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n938), .B1(KEYINPUT122), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n941), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n933), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G301), .B1(new_n931), .B2(new_n925), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n916), .A2(new_n925), .A3(G301), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n899), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT124), .B(new_n899), .C1(new_n954), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n962));
  NOR2_X1   g537(.A1(G166), .A2(new_n938), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT55), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n904), .A2(new_n914), .A3(new_n906), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n672), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n920), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT109), .B1(new_n902), .B2(new_n903), .ZN(new_n970));
  NOR3_X1   g545(.A1(G164), .A2(new_n918), .A3(G1384), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n914), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  NOR2_X1   g549(.A1(G164), .A2(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G2090), .B1(new_n977), .B2(KEYINPUT115), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n972), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n968), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n962), .B(new_n965), .C1(new_n981), .C2(new_n938), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n920), .B1(new_n917), .B2(new_n919), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n914), .B1(new_n922), .B2(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT115), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n985), .A3(new_n754), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n938), .B1(new_n986), .B2(new_n967), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT116), .B1(new_n987), .B2(new_n964), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n967), .B1(new_n924), .B2(G2090), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G8), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n964), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n996));
  OAI21_X1  g571(.A(G1981), .B1(new_n564), .B2(new_n567), .ZN(new_n997));
  INV_X1    g572(.A(G61), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n504), .B2(new_n505), .ZN(new_n999));
  INV_X1    g574(.A(new_n566), .ZN(new_n1000));
  OAI21_X1  g575(.A(G651), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n495), .A2(G86), .A3(new_n506), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n562), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n997), .A2(KEYINPUT49), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT49), .B1(new_n997), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n917), .A2(new_n919), .A3(new_n914), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(G8), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT113), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n559), .A2(G1976), .A3(new_n560), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT112), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(new_n1008), .A3(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1012), .A2(new_n1008), .A3(G8), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n996), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1009), .B(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(KEYINPUT117), .A3(new_n1017), .A4(new_n1014), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n995), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n989), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT125), .B1(new_n961), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n989), .A2(new_n1023), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT125), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n960), .A4(new_n953), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT61), .ZN(new_n1029));
  XOR2_X1   g604(.A(G299), .B(KEYINPUT57), .Z(new_n1030));
  NAND2_X1  g605(.A1(new_n977), .A2(new_n724), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT56), .B(G2072), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n907), .A2(new_n914), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1030), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1029), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(new_n1029), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1030), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT61), .A3(new_n1034), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1008), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT58), .B(G1341), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n1046), .A2(new_n1047), .B1(G1996), .B2(new_n966), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n540), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT119), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1051), .A3(new_n540), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(KEYINPUT59), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT59), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n924), .A2(new_n750), .B1(new_n1046), .B2(new_n771), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n591), .B1(new_n1057), .B2(KEYINPUT60), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(KEYINPUT60), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1041), .A2(new_n1056), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1057), .A2(new_n583), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1034), .B1(new_n1036), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1025), .A2(new_n1028), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n995), .B1(new_n965), .B2(new_n991), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n937), .A2(G286), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1010), .A2(new_n1018), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(KEYINPUT63), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n989), .A2(new_n1023), .A3(new_n1067), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n989), .A2(new_n1023), .A3(KEYINPUT118), .A4(new_n1067), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1069), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1021), .A2(new_n1015), .A3(new_n560), .A4(new_n559), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1004), .B(KEYINPUT114), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n938), .B(new_n1046), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n995), .B2(new_n1068), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT126), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n951), .A2(new_n1082), .A3(new_n952), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1026), .A2(new_n1081), .A3(new_n1083), .A4(new_n954), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n989), .A2(new_n1023), .A3(new_n954), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n936), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n934), .A2(KEYINPUT121), .A3(new_n935), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(G168), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1089), .A2(new_n949), .B1(new_n937), .B2(new_n940), .ZN(new_n1090));
  INV_X1    g665(.A(new_n952), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1090), .A2(KEYINPUT62), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT126), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT62), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1084), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1065), .A2(new_n1076), .A3(new_n1080), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n922), .A2(new_n905), .A3(new_n914), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(G1996), .A3(new_n818), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT108), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n769), .B(new_n771), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(G1996), .B2(new_n818), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n692), .B1(new_n688), .B2(new_n689), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n690), .A2(new_n693), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1098), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n575), .B(new_n686), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1098), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1096), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1097), .B1(new_n1101), .B2(new_n735), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT46), .B1(new_n1097), .B2(G1996), .ZN(new_n1112));
  OR3_X1    g687(.A1(new_n1097), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT47), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n769), .A2(G2067), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1097), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1107), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1098), .A2(new_n686), .A3(new_n575), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT48), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1115), .B(new_n1118), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1110), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g698(.A(G319), .ZN(new_n1125));
  INV_X1    g699(.A(new_n625), .ZN(new_n1126));
  NOR4_X1   g700(.A1(G229), .A2(new_n1125), .A3(new_n1126), .A4(G227), .ZN(new_n1127));
  OAI211_X1 g701(.A(new_n839), .B(new_n1127), .C1(new_n895), .C2(new_n896), .ZN(G225));
  INV_X1    g702(.A(G225), .ZN(G308));
endmodule


