//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT96), .B(G57gat), .Z(new_n208));
  INV_X1    g007(.A(G64gat), .ZN(new_n209));
  OR3_X1    g008(.A1(new_n208), .A2(KEYINPUT97), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  OR2_X1    g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n208), .A2(new_n209), .ZN(new_n215));
  INV_X1    g014(.A(G57gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT97), .B1(new_n216), .B2(G64gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n210), .B(new_n214), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G57gat), .B(G64gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n211), .B(new_n212), .C1(new_n219), .C2(new_n213), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n207), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n222), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT98), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n227), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G155gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(G211gat), .ZN(new_n232));
  AND2_X1   g031(.A1(G231gat), .A2(G233gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n230), .B(new_n234), .Z(new_n235));
  INV_X1    g034(.A(KEYINPUT99), .ZN(new_n236));
  INV_X1    g035(.A(G99gat), .ZN(new_n237));
  INV_X1    g036(.A(G106gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(KEYINPUT8), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT7), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n241), .B(new_n243), .C1(G85gat), .C2(G92gat), .ZN(new_n244));
  XOR2_X1   g043(.A(G99gat), .B(G106gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT100), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G29gat), .ZN(new_n249));
  INV_X1    g048(.A(G36gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT14), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(G29gat), .A2(G36gat), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G43gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT15), .B1(new_n258), .B2(G50gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n258), .B2(G50gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n257), .B(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G50gat), .ZN(new_n262));
  OR3_X1    g061(.A1(new_n262), .A2(KEYINPUT93), .A3(G43gat), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT93), .B1(new_n262), .B2(G43gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n263), .B(new_n264), .C1(new_n258), .C2(G50gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT15), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT41), .ZN(new_n272));
  NAND2_X1  g071(.A1(G232gat), .A2(G233gat), .ZN(new_n273));
  OAI221_X1 g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .C1(new_n268), .C2(new_n248), .ZN(new_n274));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G134gat), .B(G162gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n272), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n276), .B(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n235), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n221), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT101), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n221), .B(new_n246), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(KEYINPUT10), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n247), .A2(KEYINPUT101), .A3(KEYINPUT10), .A4(new_n282), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G230gat), .A2(G233gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT102), .ZN(new_n294));
  XNOR2_X1  g093(.A(G120gat), .B(G148gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G176gat), .B(G204gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n291), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT103), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n291), .A2(new_n293), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G127gat), .A2(G134gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G127gat), .A2(G134gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G113gat), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n308), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT69), .B1(new_n306), .B2(new_n307), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  INV_X1    g120(.A(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT1), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n315), .A2(G120gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n313), .A2(G113gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT68), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n327), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n327), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n319), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(G162gat), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT2), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G155gat), .ZN(new_n343));
  INV_X1    g142(.A(G155gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G162gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G155gat), .B(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT78), .ZN(new_n350));
  XOR2_X1   g149(.A(G141gat), .B(G148gat), .Z(new_n351));
  NAND4_X1  g150(.A1(new_n341), .A2(new_n348), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n320), .A2(new_n326), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n309), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n314), .A2(new_n316), .A3(new_n331), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n331), .B1(new_n314), .B2(new_n316), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT70), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n327), .A2(new_n333), .A3(new_n334), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n319), .A2(new_n355), .A3(new_n352), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n365), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n365), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(KEYINPUT83), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT78), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT78), .B1(new_n343), .B2(new_n345), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G141gat), .B(G148gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n340), .B2(KEYINPUT2), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n354), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n319), .C1(new_n335), .C2(new_n336), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n364), .B1(new_n377), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n363), .B(new_n361), .C1(new_n388), .C2(new_n375), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT5), .ZN(new_n390));
  INV_X1    g189(.A(new_n308), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT1), .B1(new_n317), .B2(KEYINPUT67), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n310), .A2(new_n311), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n371), .B2(new_n372), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT81), .B1(new_n395), .B2(new_n383), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n337), .A2(new_n397), .A3(new_n359), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n363), .B1(new_n399), .B2(new_n384), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n387), .B1(new_n390), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  INV_X1    g207(.A(new_n406), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n387), .B(new_n409), .C1(new_n390), .C2(new_n400), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n407), .A2(KEYINPUT84), .A3(new_n408), .A4(new_n410), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  INV_X1    g216(.A(G169gat), .ZN(new_n418));
  INV_X1    g217(.A(G176gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT26), .ZN(new_n421));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT26), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT27), .B(G183gat), .ZN(new_n427));
  INV_X1    g226(.A(G190gat), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT28), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT28), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n417), .B(new_n426), .C1(new_n429), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT66), .ZN(new_n435));
  INV_X1    g234(.A(new_n417), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(new_n432), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n426), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT23), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n422), .A2(KEYINPUT23), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n420), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT65), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n224), .A2(new_n428), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT65), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n446), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n452), .A2(new_n450), .ZN(new_n457));
  INV_X1    g256(.A(new_n447), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT25), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n456), .A2(KEYINPUT25), .B1(new_n446), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT29), .B1(new_n443), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT76), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G211gat), .A2(G218gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT22), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT74), .ZN(new_n468));
  XNOR2_X1  g267(.A(G197gat), .B(G204gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(G211gat), .A2(G218gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT75), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n465), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n468), .A3(new_n469), .A4(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT76), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n446), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n445), .A2(new_n420), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n423), .A2(KEYINPUT23), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT24), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n417), .A2(new_n448), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n448), .B1(new_n417), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n482), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n435), .B2(new_n442), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n481), .B(new_n462), .C1(new_n494), .C2(KEYINPUT29), .ZN(new_n495));
  INV_X1    g294(.A(new_n434), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT77), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT77), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n460), .A2(new_n498), .A3(new_n434), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n499), .A3(new_n463), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n464), .A2(new_n480), .A3(new_n495), .A4(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n497), .A2(new_n499), .A3(new_n503), .A4(new_n462), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n494), .A2(new_n463), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n479), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G64gat), .B(G92gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n502), .B1(new_n501), .B2(new_n506), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI211_X1 g313(.A(new_n502), .B(new_n511), .C1(new_n501), .C2(new_n506), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n416), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G228gat), .A2(G233gat), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n477), .B2(new_n478), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n520), .A2(KEYINPUT3), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n521), .B2(new_n359), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n358), .A2(new_n503), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n480), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(KEYINPUT86), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n526));
  INV_X1    g325(.A(new_n519), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n520), .A2(KEYINPUT3), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n383), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n479), .B1(new_n358), .B2(new_n503), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n519), .B(KEYINPUT85), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n473), .A2(new_n465), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT29), .B1(new_n472), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n535), .B2(new_n472), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n357), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n359), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n534), .B1(new_n539), .B2(new_n524), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(G22gat), .ZN(new_n543));
  INV_X1    g342(.A(G22gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n532), .A2(new_n544), .A3(new_n541), .ZN(new_n545));
  XNOR2_X1  g344(.A(G78gat), .B(G106gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G50gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n543), .A2(KEYINPUT88), .A3(new_n545), .A4(new_n548), .ZN(new_n552));
  INV_X1    g351(.A(new_n548), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n544), .B1(new_n532), .B2(new_n541), .ZN(new_n554));
  AOI211_X1 g353(.A(G22gat), .B(new_n540), .C1(new_n525), .C2(new_n531), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n558), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n551), .A2(new_n552), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n518), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n434), .A2(KEYINPUT66), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n441), .B1(new_n440), .B2(new_n426), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n460), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n395), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n443), .A2(new_n337), .A3(new_n460), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G227gat), .ZN(new_n569));
  INV_X1    g368(.A(G233gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT34), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n569), .A2(new_n570), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n573), .A3(new_n567), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(KEYINPUT71), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(KEYINPUT32), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G15gat), .B(G43gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G99gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT71), .B1(new_n574), .B2(new_n575), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(KEYINPUT72), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n575), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n577), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n572), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n583), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n590), .A2(new_n577), .A3(new_n581), .A4(new_n576), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n571), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n562), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n597), .A3(new_n595), .ZN(new_n598));
  OAI211_X1 g397(.A(KEYINPUT73), .B(new_n572), .C1(new_n584), .C2(new_n588), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n596), .B1(new_n600), .B2(new_n562), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n399), .A2(new_n363), .A3(new_n384), .ZN(new_n602));
  INV_X1    g401(.A(new_n361), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT83), .B1(new_n384), .B2(KEYINPUT4), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n606), .B2(new_n385), .ZN(new_n607));
  OAI211_X1 g406(.A(KEYINPUT39), .B(new_n602), .C1(new_n607), .C2(new_n363), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n361), .B1(new_n377), .B2(new_n386), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610));
  INV_X1    g409(.A(new_n363), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n608), .A2(KEYINPUT40), .A3(new_n612), .A4(new_n409), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n613), .A2(new_n407), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n409), .A3(new_n612), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT40), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n516), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n551), .A2(new_n552), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n557), .A2(new_n559), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n411), .A2(KEYINPUT89), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n407), .A2(new_n623), .A3(new_n408), .A4(new_n410), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n414), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n501), .A2(new_n506), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT37), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT38), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n464), .A2(new_n500), .A3(new_n495), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n479), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n504), .A2(new_n505), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(KEYINPUT37), .C1(new_n479), .C2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(new_n632), .A3(new_n510), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n511), .B1(new_n626), .B2(KEYINPUT38), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n626), .B(KEYINPUT37), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n618), .B(new_n621), .C1(new_n625), .C2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n561), .A2(new_n601), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT35), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n600), .A2(new_n621), .A3(new_n517), .A4(new_n625), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n589), .A2(new_n595), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n560), .A2(new_n642), .A3(new_n640), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n416), .A2(new_n517), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n640), .A2(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n305), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n268), .A2(new_n207), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n270), .B2(new_n207), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT18), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT94), .B1(new_n268), .B2(new_n207), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n647), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n649), .B(KEYINPUT13), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT91), .ZN(new_n658));
  XOR2_X1   g457(.A(G169gat), .B(G197gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n651), .A2(new_n655), .A3(new_n656), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT95), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n666));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n665), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n416), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n671), .A2(new_n517), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(KEYINPUT42), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n206), .B2(new_n678), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n671), .A2(new_n685), .A3(new_n601), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n672), .A2(new_n600), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n671), .A2(new_n621), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NAND2_X1  g490(.A1(new_n639), .A2(KEYINPUT108), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n561), .A2(new_n601), .A3(new_n638), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n645), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n695), .B2(new_n280), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  INV_X1    g496(.A(new_n280), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n697), .B(new_n698), .C1(new_n645), .C2(new_n639), .ZN(new_n699));
  INV_X1    g498(.A(new_n235), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n669), .A2(new_n700), .A3(new_n303), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n416), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n698), .B1(new_n645), .B2(new_n639), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n701), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(G29gat), .A3(new_n416), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n710), .ZN(G1328gat));
  OAI21_X1  g510(.A(G36gat), .B1(new_n704), .B2(new_n517), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n707), .A2(G36gat), .A3(new_n517), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT46), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(G1329gat));
  NAND4_X1  g514(.A1(new_n706), .A2(new_n258), .A3(new_n600), .A4(new_n701), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n696), .A2(new_n601), .A3(new_n699), .A4(new_n702), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n258), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n720), .B(new_n716), .C1(new_n717), .C2(new_n258), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT47), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(new_n262), .B1(new_n707), .B2(new_n621), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n560), .A2(G50gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n704), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g527(.A1(new_n695), .A2(new_n281), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n670), .A2(new_n304), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n416), .B(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n208), .ZN(G1332gat));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n517), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n731), .A2(new_n742), .A3(new_n600), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  OAI21_X1  g543(.A(G71gat), .B1(new_n735), .B2(new_n601), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n748), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(KEYINPUT50), .A3(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n560), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n696), .A2(new_n699), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n670), .A2(new_n700), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n303), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G85gat), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n757), .A2(new_n758), .A3(new_n416), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n695), .A2(KEYINPUT51), .A3(new_n280), .A4(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n695), .A2(new_n280), .A3(new_n756), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n695), .A2(new_n280), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n769), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n756), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(KEYINPUT113), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n765), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(new_n673), .A3(new_n303), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n759), .B1(new_n774), .B2(new_n758), .ZN(G1336gat));
  NOR2_X1   g574(.A1(new_n517), .A2(G92gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n303), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n516), .A3(new_n303), .A4(new_n756), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(new_n778), .B2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n766), .A2(KEYINPUT115), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n766), .B2(new_n781), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n761), .B(KEYINPUT112), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n303), .B(new_n776), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n778), .A2(G92gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n780), .A2(new_n789), .ZN(G1337gat));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n757), .A2(new_n791), .A3(new_n601), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n757), .B2(new_n601), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(G99gat), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n773), .A2(new_n237), .A3(new_n600), .A4(new_n303), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1338gat));
  NOR3_X1   g595(.A1(new_n304), .A2(G106gat), .A3(new_n621), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n773), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n755), .A2(new_n560), .A3(new_n303), .A4(new_n756), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n238), .A2(KEYINPUT117), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n238), .A2(KEYINPUT117), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n797), .ZN(new_n805));
  INV_X1    g604(.A(new_n784), .ZN(new_n806));
  INV_X1    g605(.A(new_n785), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n803), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT53), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n810), .ZN(G1339gat));
  NOR2_X1   g610(.A1(new_n653), .A2(new_n654), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n648), .A2(new_n649), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n662), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n664), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n280), .B1(new_n303), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n285), .A2(new_n292), .A3(new_n287), .A4(new_n288), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n291), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT118), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n291), .A2(new_n820), .A3(KEYINPUT54), .A4(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n291), .A2(KEYINPUT54), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n298), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n300), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n816), .B1(new_n669), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n827), .A2(new_n300), .A3(new_n828), .A4(new_n815), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n700), .B1(new_n831), .B2(new_n280), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n235), .A2(new_n280), .A3(new_n303), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n669), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n732), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n560), .A2(new_n642), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n837), .A2(new_n517), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n670), .A2(new_n315), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT119), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n416), .A2(new_n516), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n836), .A2(new_n621), .A3(new_n600), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n669), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(G1340gat));
  NAND3_X1  g645(.A1(new_n839), .A2(new_n313), .A3(new_n303), .ZN(new_n847));
  OAI21_X1  g646(.A(G120gat), .B1(new_n844), .B2(new_n304), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1341gat));
  NOR3_X1   g648(.A1(new_n844), .A2(new_n321), .A3(new_n235), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n839), .A2(new_n700), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n321), .ZN(G1342gat));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n517), .A3(new_n838), .A4(new_n280), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT56), .B1(new_n853), .B2(G134gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n853), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(KEYINPUT56), .C1(new_n853), .C2(G134gat), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n844), .B2(new_n698), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n855), .A2(new_n856), .A3(new_n858), .A4(new_n859), .ZN(G1343gat));
  INV_X1    g659(.A(G141gat), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n601), .A2(new_n560), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n837), .A2(new_n517), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n669), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n836), .A2(new_n865), .A3(new_n560), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n830), .A2(new_n832), .B1(new_n669), .B2(new_n834), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT57), .B1(new_n867), .B2(new_n621), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n866), .A2(new_n868), .A3(new_n601), .A4(new_n843), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n670), .A2(G141gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n864), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n864), .B(KEYINPUT58), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1344gat));
  OR3_X1    g674(.A1(new_n863), .A2(G148gat), .A3(new_n304), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  INV_X1    g676(.A(new_n869), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n303), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n877), .B(G148gat), .C1(new_n869), .C2(new_n304), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n876), .B1(new_n880), .B2(new_n882), .ZN(G1345gat));
  INV_X1    g682(.A(new_n863), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n884), .A2(new_n700), .B1(new_n338), .B2(new_n339), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n700), .A2(new_n338), .A3(new_n339), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n878), .B2(new_n886), .ZN(G1346gat));
  OR3_X1    g686(.A1(new_n869), .A2(KEYINPUT121), .A3(new_n698), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT121), .B1(new_n869), .B2(new_n698), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(G162gat), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n342), .A3(new_n280), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n867), .A2(new_n673), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(new_n516), .A3(new_n838), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n418), .A3(new_n670), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n732), .A2(new_n517), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n600), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(KEYINPUT122), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n621), .B1(new_n897), .B2(KEYINPUT122), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n867), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n669), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n895), .A2(new_n901), .ZN(G1348gat));
  NAND3_X1  g701(.A1(new_n894), .A2(new_n419), .A3(new_n303), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  OAI21_X1  g703(.A(G176gat), .B1(new_n900), .B2(new_n304), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n894), .A2(new_n427), .A3(new_n700), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n900), .A2(new_n235), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n224), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n909), .B(new_n913), .C1(new_n224), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1350gat));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n428), .A3(new_n280), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n900), .A2(new_n698), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n917), .A2(new_n918), .A3(G190gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n917), .B2(G190gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(G1351gat));
  NAND4_X1  g720(.A1(new_n866), .A2(new_n868), .A3(new_n601), .A4(new_n896), .ZN(new_n922));
  OR3_X1    g721(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n669), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT124), .B1(new_n922), .B2(new_n669), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(G197gat), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n893), .A2(new_n516), .A3(new_n862), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n670), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(G1352gat));
  INV_X1    g728(.A(new_n922), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(KEYINPUT125), .A3(new_n303), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n922), .B2(new_n304), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(G204gat), .A3(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n926), .A2(new_n935), .A3(new_n303), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(G1353gat));
  INV_X1    g738(.A(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n930), .B2(new_n700), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(KEYINPUT63), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT63), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n940), .A3(new_n700), .ZN(new_n946));
  OAI21_X1  g745(.A(G211gat), .B1(new_n922), .B2(new_n235), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n942), .A3(KEYINPUT63), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n926), .B2(new_n280), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n280), .A2(G218gat), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT127), .Z(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n930), .B2(new_n952), .ZN(G1355gat));
endmodule


