//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n461), .B1(new_n455), .B2(new_n451), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n471), .B(G125), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(G137), .B(new_n478), .C1(new_n473), .C2(new_n474), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n468), .A2(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G137), .A4(new_n478), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n467), .A2(G2105), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n480), .A2(new_n483), .B1(G101), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n477), .A2(new_n485), .ZN(G160));
  AOI21_X1  g061(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n478), .B1(new_n468), .B2(new_n469), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NOR2_X1   g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(new_n478), .B2(G112), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n488), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT71), .ZN(G162));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n473), .B2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT72), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(new_n495), .C1(new_n473), .C2(new_n474), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT4), .A2(G138), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n467), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n487), .A2(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n478), .C1(new_n473), .C2(new_n474), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n500), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT73), .B(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n513), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n515), .A2(G50), .B1(G75), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(new_n522), .A3(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(new_n522), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n519), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n515), .A2(G51), .A3(G543), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n515), .A2(G89), .A3(new_n522), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n520), .A2(new_n521), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n547), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n516), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n515), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n524), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT76), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n546), .A2(new_n516), .A3(new_n548), .ZN(new_n555));
  INV_X1    g130(.A(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n514), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n511), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n518), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G52), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n561), .A2(new_n543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G90), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n555), .A2(new_n563), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n554), .A2(new_n567), .ZN(G171));
  NAND2_X1  g143(.A1(new_n564), .A2(G81), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n562), .A2(G43), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n513), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  NAND4_X1  g150(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  NAND2_X1  g155(.A1(new_n522), .A2(G65), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT80), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n556), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g159(.A(G91), .B(new_n522), .C1(new_n560), .C2(new_n511), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT79), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n515), .A2(new_n587), .A3(G91), .A4(new_n522), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT9), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(G53), .B(G543), .C1(new_n560), .C2(new_n511), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT78), .B(KEYINPUT9), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n589), .A2(new_n596), .ZN(G299));
  INV_X1    g172(.A(G171), .ZN(G301));
  NAND2_X1  g173(.A1(new_n540), .A2(KEYINPUT81), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n537), .A2(new_n538), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n600), .A2(new_n601), .A3(new_n539), .A4(new_n536), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G286));
  NAND3_X1  g179(.A1(new_n515), .A2(G87), .A3(new_n522), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n515), .A2(G49), .A3(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G288));
  NAND3_X1  g183(.A1(new_n515), .A2(G86), .A3(new_n522), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n515), .A2(G48), .A3(G543), .ZN(new_n610));
  INV_X1    g185(.A(G61), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n520), .B2(new_n521), .ZN(new_n612));
  AND2_X1   g187(.A1(G73), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n516), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(G305));
  INV_X1    g190(.A(G47), .ZN(new_n616));
  INV_X1    g191(.A(G85), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n616), .A2(new_n551), .B1(new_n524), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT82), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(new_n513), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(G290));
  INV_X1    g197(.A(G54), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n522), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n624));
  OAI22_X1  g199(.A1(new_n551), .A2(new_n623), .B1(new_n556), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n564), .A2(KEYINPUT10), .A3(G92), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n524), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G868), .B2(G171), .ZN(G284));
  XNOR2_X1  g208(.A(G284), .B(KEYINPUT83), .ZN(G321));
  NOR2_X1   g209(.A1(G299), .A2(G868), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n603), .ZN(G297));
  AOI21_X1  g211(.A(new_n635), .B1(G868), .B2(new_n603), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n630), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n630), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n574), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n489), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(new_n478), .B2(G111), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n487), .A2(KEYINPUT85), .A3(G135), .ZN(new_n647));
  AOI21_X1  g222(.A(KEYINPUT85), .B1(new_n487), .B2(G135), .ZN(new_n648));
  OAI221_X1 g223(.A(new_n644), .B1(new_n645), .B2(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n481), .A2(new_n484), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT84), .B(G2100), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(G2096), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n655), .B(new_n656), .C1(new_n653), .C2(new_n654), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT86), .Z(G156));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT87), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2438), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2427), .B(G2430), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n666), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n669), .ZN(new_n673));
  OAI21_X1  g248(.A(G14), .B1(new_n665), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(new_n665), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT89), .ZN(G401));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT17), .Z(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(new_n677), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n682), .C1(new_n680), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n677), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1971), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n695), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n701), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1981), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n706), .B1(new_n701), .B2(new_n705), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n693), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n714), .A2(new_n692), .A3(new_n710), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(G1991), .B(G1996), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT92), .B(G1986), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n718), .A2(new_n722), .A3(new_n720), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(G229));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G32), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT26), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G129), .B2(new_n489), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n487), .A2(G141), .B1(G105), .B2(new_n484), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT103), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT27), .B(G1996), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n630), .B2(new_n739), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1348), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n727), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n727), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(G2078), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G28), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT104), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n749), .B(new_n727), .C1(new_n747), .C2(G28), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n746), .B(new_n750), .C1(new_n649), .C2(new_n727), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n727), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n487), .A2(G139), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n481), .A2(G127), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n478), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n752), .B1(new_n760), .B2(new_n727), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n751), .B1(new_n761), .B2(G2072), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G2078), .B2(new_n744), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n738), .A2(new_n742), .A3(new_n745), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n739), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n574), .B2(new_n739), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT97), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1341), .ZN(new_n768));
  NOR2_X1   g343(.A1(G5), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G171), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n764), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n761), .A2(G2072), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT102), .Z(new_n775));
  NOR2_X1   g350(.A1(G160), .A2(new_n727), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n727), .B1(KEYINPUT24), .B2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(KEYINPUT24), .B2(G34), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n727), .A2(G26), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT100), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n487), .A2(G140), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT98), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n788));
  INV_X1    g363(.A(G104), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n478), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n489), .A2(G128), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n489), .A2(KEYINPUT99), .A3(G128), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n785), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT101), .B(G2067), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n775), .A2(new_n781), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n727), .A2(G35), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT105), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n727), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT29), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G2090), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n739), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n739), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n780), .B2(new_n779), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n801), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n805), .A2(G2090), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n739), .A2(G20), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT23), .Z(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G299), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1956), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT106), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n773), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n739), .A2(G24), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT93), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n619), .A2(new_n621), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n739), .ZN(new_n824));
  INV_X1    g399(.A(G1986), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n727), .A2(G25), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n489), .A2(G119), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n487), .A2(G131), .ZN(new_n829));
  OR2_X1    g404(.A1(G95), .A2(G2105), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n827), .B1(new_n833), .B2(new_n727), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT35), .B(G1991), .Z(new_n835));
  XOR2_X1   g410(.A(new_n834), .B(new_n835), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(G303), .A2(G16), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n739), .A2(G22), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT94), .B(G1971), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n847));
  MUX2_X1   g422(.A(G23), .B(G288), .S(G16), .Z(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT33), .B(G1976), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  MUX2_X1   g425(.A(G6), .B(G305), .S(G16), .Z(new_n851));
  XOR2_X1   g426(.A(KEYINPUT32), .B(G1981), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n846), .A2(new_n847), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n844), .A3(new_n845), .ZN(new_n855));
  INV_X1    g430(.A(new_n850), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT95), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT34), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n838), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT34), .B1(new_n854), .B2(new_n857), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n826), .A2(new_n837), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT96), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n858), .A2(new_n859), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT36), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT36), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n820), .B1(new_n870), .B2(new_n872), .ZN(G311));
  INV_X1    g448(.A(new_n820), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n871), .B1(new_n866), .B2(new_n868), .ZN(new_n875));
  AOI211_X1 g450(.A(KEYINPUT36), .B(new_n867), .C1(new_n862), .C2(new_n865), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(G150));
  XOR2_X1   g452(.A(KEYINPUT107), .B(G55), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n562), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n564), .A2(G93), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(new_n513), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n883), .A2(new_n573), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n573), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT38), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n631), .A2(new_n638), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n890));
  AOI21_X1  g465(.A(G860), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n890), .B2(new_n889), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n883), .A2(G860), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT37), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(G145));
  XNOR2_X1  g470(.A(G162), .B(new_n649), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G160), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n733), .B(new_n832), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n796), .B(G164), .ZN(new_n900));
  INV_X1    g475(.A(new_n760), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n652), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n489), .A2(G130), .ZN(new_n905));
  NOR2_X1   g480(.A1(G106), .A2(G2105), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(new_n478), .B2(G118), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n487), .A2(KEYINPUT108), .A3(G142), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT108), .B1(new_n487), .B2(G142), .ZN(new_n909));
  OAI221_X1 g484(.A(new_n905), .B1(new_n906), .B2(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n652), .A3(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n900), .A2(new_n901), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n903), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n903), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n899), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n918), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n914), .B(new_n916), .C1(new_n922), .C2(new_n902), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n903), .A2(new_n917), .A3(new_n918), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n898), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n897), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n921), .A2(new_n897), .A3(new_n925), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g508(.A(G290), .B(G305), .ZN(new_n934));
  XNOR2_X1  g509(.A(G303), .B(G288), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n934), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n823), .A2(G305), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n823), .A2(G305), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n934), .A2(new_n935), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT42), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n883), .B(new_n573), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(new_n640), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n630), .A2(G299), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n630), .A2(G299), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n948), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT41), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n948), .B(KEYINPUT111), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n951), .A2(KEYINPUT41), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n960), .A2(new_n947), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n938), .A2(new_n945), .A3(new_n953), .A4(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n953), .B1(new_n960), .B2(new_n947), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(new_n943), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n963), .B1(new_n966), .B2(new_n944), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G868), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  INV_X1    g545(.A(G868), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n883), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n962), .B2(new_n967), .ZN(new_n974));
  INV_X1    g549(.A(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT112), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(G295));
  NAND2_X1  g552(.A1(new_n969), .A2(new_n972), .ZN(G331));
  AND3_X1   g553(.A1(new_n554), .A2(new_n540), .A3(new_n567), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n554), .A2(new_n567), .B1(new_n602), .B2(new_n599), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n946), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G171), .A2(new_n603), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n554), .A2(new_n540), .A3(new_n567), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n886), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(KEYINPUT113), .B(new_n946), .C1(new_n979), .C2(new_n980), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n986), .A2(new_n959), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n951), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n957), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n981), .A2(new_n984), .A3(KEYINPUT114), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n946), .C1(new_n979), .C2(new_n980), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n937), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n993), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n952), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n986), .A2(new_n959), .A3(new_n987), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n964), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G37), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n958), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n952), .A2(new_n955), .B1(new_n948), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(new_n996), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n990), .B1(new_n986), .B2(new_n987), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n937), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND4_X1   g583(.A1(KEYINPUT43), .A2(new_n1008), .A3(new_n1000), .A4(new_n999), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT44), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1008), .A2(new_n1002), .A3(new_n1000), .A4(new_n999), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(G397));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n487), .A2(new_n501), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n504), .A2(new_n502), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n508), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n498), .B1(new_n481), .B2(new_n495), .ZN(new_n1023));
  INV_X1    g598(.A(new_n499), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1019), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n477), .A2(G40), .A3(new_n485), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n509), .A2(new_n1031), .A3(new_n1019), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(G2090), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G1384), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n509), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1026), .A2(new_n1036), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n509), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1030), .ZN(new_n1042));
  INV_X1    g617(.A(G1971), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1018), .B1(new_n1034), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1017), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n509), .A2(new_n1019), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1030), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n605), .A2(new_n606), .A3(G1976), .A4(new_n607), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(G8), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n477), .A2(new_n485), .A3(G40), .ZN(new_n1056));
  OAI211_X1 g631(.A(G8), .B(new_n1052), .C1(new_n1056), .C2(new_n1026), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT52), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n609), .A2(new_n610), .A3(new_n708), .A4(new_n614), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(KEYINPUT49), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1051), .A3(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT49), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1055), .B(new_n1058), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n509), .A2(new_n1019), .A3(new_n1027), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1030), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1018), .B1(new_n1044), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1064), .B1(new_n1069), .B2(new_n1048), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1041), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(new_n1038), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT45), .B1(new_n509), .B2(new_n1019), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n1056), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1971), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1033), .A2(G2090), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1046), .B(KEYINPUT55), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(KEYINPUT119), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n509), .A2(new_n1037), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n809), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1065), .A2(new_n1030), .A3(new_n780), .A4(new_n1067), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1018), .B(G286), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1049), .A2(new_n1070), .A3(new_n1079), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT120), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1069), .A2(new_n1048), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1091), .A2(new_n1070), .A3(KEYINPUT63), .A4(new_n1084), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1060), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G288), .A2(G1976), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1051), .A2(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1069), .A2(new_n1048), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1097), .A2(new_n1098), .B1(new_n1099), .B2(new_n1064), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1040), .A2(new_n1080), .A3(new_n1030), .ZN(new_n1102));
  OAI211_X1 g677(.A(G168), .B(new_n1083), .C1(new_n1102), .C2(G1966), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(G168), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT51), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1107), .A3(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1101), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1049), .A2(new_n1070), .A3(new_n1079), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1042), .B2(G2078), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1102), .A2(KEYINPUT53), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1065), .A2(new_n1030), .A3(new_n1067), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n771), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G171), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1109), .A2(new_n1110), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1106), .A2(new_n1101), .A3(new_n1108), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1100), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n596), .B2(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G299), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n589), .B(new_n596), .C1(KEYINPUT122), .C2(KEYINPUT57), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1074), .A2(new_n1039), .A3(new_n1041), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT121), .B(G1956), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1033), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT123), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1125), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G1348), .ZN(new_n1138));
  INV_X1    g713(.A(G2067), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1056), .A2(new_n1026), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1115), .A2(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n631), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1134), .A2(new_n1142), .A3(KEYINPUT124), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(KEYINPUT125), .ZN(new_n1149));
  INV_X1    g724(.A(G1996), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1074), .A2(new_n1150), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1051), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1149), .B1(new_n1154), .B2(new_n574), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1149), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n573), .B(new_n1156), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n631), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1115), .A2(new_n1138), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1051), .A2(G2067), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n630), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1158), .A2(new_n1159), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1170), .B2(KEYINPUT126), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1172), .A3(new_n1169), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1147), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1050), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT45), .B1(new_n1026), .B2(KEYINPUT115), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1056), .A2(new_n1111), .A3(G2078), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1072), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1112), .A2(new_n1180), .A3(new_n1116), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(G171), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1112), .A2(new_n1114), .A3(G301), .A4(new_n1116), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1182), .A2(KEYINPUT54), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1184), .A2(new_n1110), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1112), .A2(new_n1180), .A3(G301), .A4(new_n1116), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT54), .B1(new_n1118), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g765(.A(KEYINPUT127), .B(KEYINPUT54), .C1(new_n1118), .C2(new_n1187), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1185), .B(new_n1186), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1093), .B(new_n1121), .C1(new_n1174), .C2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1178), .A2(new_n1056), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n796), .B(new_n1139), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n733), .B(new_n1150), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n832), .B(new_n835), .Z(new_n1198));
  OAI21_X1  g773(.A(new_n1194), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(G290), .B(new_n825), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1194), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT116), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1193), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n833), .A2(new_n835), .ZN(new_n1205));
  OAI22_X1  g780(.A1(new_n1197), .A2(new_n1205), .B1(G2067), .B2(new_n796), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1194), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n823), .A2(new_n1194), .A3(new_n825), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1199), .B1(new_n1209), .B2(KEYINPUT48), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT48), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1194), .A2(new_n1150), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT46), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1195), .A2(new_n734), .ZN(new_n1215));
  AOI22_X1  g790(.A1(new_n1213), .A2(new_n1214), .B1(new_n1215), .B2(new_n1194), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1216), .B1(new_n1214), .B2(new_n1213), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT47), .ZN(new_n1218));
  OAI221_X1 g793(.A(new_n1207), .B1(new_n1210), .B2(new_n1212), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1219), .B1(new_n1218), .B2(new_n1217), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1204), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g796(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n1223), .B1(new_n724), .B2(new_n725), .ZN(new_n1224));
  NAND3_X1  g798(.A1(new_n1224), .A2(new_n1013), .A3(new_n932), .ZN(G225));
  INV_X1    g799(.A(G225), .ZN(G308));
endmodule


