//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G43gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G99gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G113gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G120gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(KEYINPUT72), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT72), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n214), .B1(new_n210), .B2(new_n211), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n209), .A2(G113gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G127gat), .A2(G134gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G127gat), .A2(G134gat), .ZN(new_n223));
  OR2_X1    g022(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g023(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n216), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n214), .A2(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n219), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n222), .ZN(new_n232));
  OR2_X1    g031(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(G134gat), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n228), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n209), .A2(G113gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n221), .B1(new_n239), .B2(new_n229), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(KEYINPUT70), .A3(new_n235), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n227), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  INV_X1    g048(.A(G176gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n245), .A2(new_n246), .A3(new_n247), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT68), .B1(new_n252), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n256));
  AND2_X1   g055(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n257));
  AND2_X1   g056(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT28), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT27), .B(G183gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n254), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(G183gat), .B1(new_n262), .B2(new_n263), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n249), .A2(new_n250), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n270), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n278));
  INV_X1    g077(.A(new_n276), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n247), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT25), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n247), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(new_n286), .B2(new_n276), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT64), .B(G169gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n275), .A2(G176gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT25), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n272), .B(new_n273), .C1(G183gat), .C2(G190gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n242), .B1(new_n269), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n276), .A2(new_n275), .ZN(new_n296));
  AND3_X1   g095(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n257), .B2(new_n256), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n296), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n295), .B1(new_n302), .B2(new_n287), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n252), .A2(new_n253), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n253), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n266), .B1(new_n264), .B2(new_n265), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  AND4_X1   g112(.A1(KEYINPUT70), .A2(new_n231), .A3(new_n222), .A4(new_n235), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT70), .B1(new_n240), .B2(new_n235), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n305), .A2(new_n313), .A3(new_n227), .A4(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n207), .B1(new_n294), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n206), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n207), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n269), .A2(new_n242), .A3(new_n293), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n305), .A2(new_n313), .B1(new_n316), .B2(new_n227), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT74), .B1(new_n318), .B2(KEYINPUT33), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n206), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n318), .A2(new_n319), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n203), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n324), .B2(KEYINPUT32), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n318), .A2(KEYINPUT74), .A3(KEYINPUT33), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n332), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT75), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n322), .A2(new_n323), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n207), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT34), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT34), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n343), .A3(new_n207), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n333), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n347));
  INV_X1    g146(.A(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(G211gat), .A2(G218gat), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G211gat), .ZN(new_n359));
  INV_X1    g158(.A(G218gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT78), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n371), .B(new_n372), .C1(new_n366), .C2(new_n365), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n364), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G197gat), .ZN(new_n375));
  INV_X1    g174(.A(G204gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n368), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n379), .A2(new_n358), .A3(new_n372), .A4(new_n363), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  INV_X1    g181(.A(G155gat), .ZN(new_n383));
  INV_X1    g182(.A(G162gat), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT82), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT82), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G148gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G141gat), .ZN(new_n390));
  INV_X1    g189(.A(G141gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G148gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n394));
  NAND2_X1  g193(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n382), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G155gat), .A2(G162gat), .ZN(new_n399));
  AND2_X1   g198(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n400));
  NOR2_X1   g199(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n397), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n388), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  OR3_X1    g205(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n406), .A2(new_n393), .B1(new_n407), .B2(new_n399), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT85), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n404), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n381), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT84), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n402), .A3(new_n393), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n416), .A2(new_n388), .B1(new_n408), .B2(new_n409), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT77), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n362), .B1(new_n361), .B2(new_n355), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n373), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n379), .A2(new_n372), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n412), .B(new_n380), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n405), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(G22gat), .B1(new_n413), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n405), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n404), .A2(new_n410), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G22gat), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n417), .B2(new_n405), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n427), .B(new_n428), .C1(new_n429), .C2(new_n381), .ZN(new_n430));
  INV_X1    g229(.A(G228gat), .ZN(new_n431));
  INV_X1    g230(.A(G233gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n424), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n424), .B2(new_n430), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n354), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n374), .A2(new_n380), .ZN(new_n438));
  INV_X1    g237(.A(new_n387), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n399), .B1(new_n439), .B2(new_n385), .ZN(new_n440));
  XNOR2_X1  g239(.A(G141gat), .B(G148gat), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n414), .B2(KEYINPUT84), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(new_n402), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n391), .A2(G148gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n389), .A2(G141gat), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n406), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n407), .A2(new_n399), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n446), .A2(new_n447), .A3(new_n409), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n443), .A2(KEYINPUT3), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n438), .B1(new_n449), .B2(KEYINPUT29), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n428), .B1(new_n450), .B2(new_n427), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n413), .A2(new_n423), .A3(G22gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n433), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n424), .A2(new_n430), .A3(new_n434), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n351), .B(KEYINPUT89), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n327), .A2(new_n328), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n332), .B1(new_n458), .B2(new_n334), .ZN(new_n459));
  INV_X1    g258(.A(new_n345), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n346), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n346), .B2(new_n461), .ZN(new_n464));
  XOR2_X1   g263(.A(G57gat), .B(G85gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n426), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n242), .A3(new_n411), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT4), .B1(new_n242), .B2(new_n426), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT4), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n316), .A2(new_n417), .A3(new_n478), .A4(new_n227), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n476), .B2(new_n479), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n472), .B(new_n475), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n479), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n473), .A3(new_n472), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n242), .A2(new_n426), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n316), .A2(new_n417), .A3(new_n227), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n474), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(KEYINPUT5), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n470), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n489), .A3(new_n470), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n490), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n497));
  AND2_X1   g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n305), .A2(new_n313), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(KEYINPUT29), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n305), .B2(new_n313), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n381), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n500), .B1(new_n269), .B2(new_n293), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n305), .A2(new_n313), .A3(new_n498), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n438), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n504), .A2(KEYINPUT79), .A3(new_n505), .A4(new_n438), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G8gat), .B(G36gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G64gat), .B(G92gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n497), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT81), .B(new_n513), .C1(new_n508), .C2(new_n509), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n496), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n508), .A2(KEYINPUT80), .A3(new_n509), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n495), .A2(new_n517), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n463), .A2(new_n464), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n202), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n346), .A2(new_n461), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n528));
  AND4_X1   g327(.A1(new_n495), .A2(new_n517), .A3(new_n521), .A4(new_n522), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n346), .A2(new_n461), .A3(new_n462), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n490), .B(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n492), .A2(new_n493), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n490), .A2(KEYINPUT92), .A3(KEYINPUT6), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT92), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n521), .A3(new_n522), .ZN(new_n541));
  INV_X1    g340(.A(new_n457), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n525), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OR3_X1    g343(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT76), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n459), .A2(new_n460), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n345), .B1(new_n329), .B2(new_n332), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT76), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n540), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n526), .A2(new_n532), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n519), .A2(KEYINPUT37), .A3(new_n520), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n514), .B1(new_n510), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT38), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n515), .ZN(new_n558));
  INV_X1    g357(.A(new_n516), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n503), .A2(new_n506), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT38), .B1(new_n560), .B2(KEYINPUT37), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n558), .A2(new_n559), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n536), .A2(new_n557), .A3(new_n539), .A4(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT39), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(new_n474), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n564), .A2(new_n474), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT39), .B1(new_n487), .B2(new_n474), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT90), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n470), .B(new_n566), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n541), .A2(new_n572), .A3(new_n534), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n563), .A2(new_n574), .A3(new_n542), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n346), .A2(KEYINPUT36), .A3(new_n546), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n549), .B2(KEYINPUT36), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n523), .A2(new_n457), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n552), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G15gat), .B(G22gat), .ZN(new_n581));
  INV_X1    g380(.A(G1gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT16), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(G1gat), .B2(new_n581), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G8gat), .ZN(new_n586));
  XOR2_X1   g385(.A(G57gat), .B(G64gat), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  INV_X1    g388(.A(G71gat), .ZN(new_n590));
  INV_X1    g389(.A(G78gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G71gat), .B(G78gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n586), .B1(KEYINPUT21), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT101), .ZN(new_n597));
  AND2_X1   g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n595), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n599), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G43gat), .B(G50gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT15), .ZN(new_n613));
  NAND2_X1  g412(.A1(G29gat), .A2(G36gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(G29gat), .A2(G36gat), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT14), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(KEYINPUT15), .B2(new_n612), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT96), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n614), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT95), .B1(new_n618), .B2(new_n619), .ZN(new_n626));
  OAI211_X1 g425(.A(KEYINPUT15), .B(new_n612), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n615), .B2(new_n621), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n623), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(G92gat), .ZN(new_n634));
  INV_X1    g433(.A(G85gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(KEYINPUT8), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G99gat), .B(G106gat), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n644), .A2(new_n636), .A3(new_n637), .A4(new_n640), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n641), .B2(new_n642), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OR3_X1    g448(.A1(new_n632), .A2(new_n633), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n649), .A2(new_n630), .B1(KEYINPUT41), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G134gat), .B(G162gat), .Z(new_n654));
  AND2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n651), .A2(KEYINPUT41), .ZN(new_n658));
  XNOR2_X1  g457(.A(G190gat), .B(G218gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n655), .B2(new_n656), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n643), .A2(new_n645), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n647), .ZN(new_n667));
  INV_X1    g466(.A(new_n648), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n600), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n595), .A2(new_n666), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT10), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  NOR4_X1   g471(.A1(new_n600), .A2(new_n646), .A3(new_n672), .A4(new_n648), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n665), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n665), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(new_n675), .A3(new_n670), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n674), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n611), .A2(new_n664), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n586), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n630), .B2(new_n631), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n632), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(G229gat), .A2(G233gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n630), .A2(new_n586), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n688), .A2(KEYINPUT18), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n689), .B(new_n690), .C1(new_n632), .C2(new_n687), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT18), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n630), .A2(KEYINPUT97), .A3(new_n586), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT97), .B1(new_n630), .B2(new_n586), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n690), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n689), .B(KEYINPUT13), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n691), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(G113gat), .B(G141gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n375), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT11), .B(G169gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT12), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n692), .A2(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n708), .B2(new_n691), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT98), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n700), .A2(new_n706), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n708), .A2(new_n691), .A3(new_n705), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n685), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n580), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n495), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT104), .B(G1gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1324gat));
  INV_X1    g519(.A(new_n541), .ZN(new_n721));
  OAI21_X1  g520(.A(G8gat), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT42), .ZN(new_n723));
  AND2_X1   g522(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n717), .A2(new_n721), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  MUX2_X1   g525(.A(new_n723), .B(KEYINPUT42), .S(new_n726), .Z(G1325gat));
  INV_X1    g526(.A(new_n717), .ZN(new_n728));
  INV_X1    g527(.A(new_n577), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n728), .A2(G15gat), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(G15gat), .B1(new_n728), .B2(new_n549), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1326gat));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n542), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(new_n664), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n609), .A2(new_n610), .ZN(new_n738));
  INV_X1    g537(.A(new_n715), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n684), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n495), .ZN(new_n742));
  INV_X1    g541(.A(G29gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n580), .A2(new_n737), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT45), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n707), .A2(new_n709), .ZN(new_n749));
  INV_X1    g548(.A(new_n684), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n611), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT105), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n550), .B1(new_n754), .B2(new_n202), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(new_n532), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT44), .B1(new_n756), .B2(new_n664), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n580), .A2(new_n758), .A3(new_n737), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n752), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n743), .B1(new_n760), .B2(new_n742), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n736), .B1(new_n748), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n758), .B1(new_n580), .B2(new_n737), .ZN(new_n763));
  AOI211_X1 g562(.A(KEYINPUT44), .B(new_n664), .C1(new_n552), .C2(new_n579), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n765), .A2(new_n495), .A3(new_n752), .ZN(new_n766));
  OAI211_X1 g565(.A(KEYINPUT106), .B(new_n747), .C1(new_n766), .C2(new_n743), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n767), .ZN(G1328gat));
  NOR2_X1   g567(.A1(new_n756), .A2(new_n664), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n741), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n770), .A2(G36gat), .A3(new_n721), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n760), .A2(new_n541), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G36gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1329gat));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n776));
  INV_X1    g575(.A(G43gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n549), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g577(.A1(new_n756), .A2(new_n664), .A3(new_n740), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n752), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n729), .B(new_n780), .C1(new_n763), .C2(new_n764), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(G43gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n777), .B1(new_n760), .B2(new_n729), .ZN(new_n785));
  OAI211_X1 g584(.A(KEYINPUT107), .B(KEYINPUT47), .C1(new_n785), .C2(new_n779), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n784), .A2(new_n786), .ZN(G1330gat));
  AOI21_X1  g586(.A(new_n348), .B1(new_n760), .B2(new_n457), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n770), .A2(G50gat), .A3(new_n542), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1331gat));
  INV_X1    g592(.A(new_n749), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n738), .A2(new_n794), .A3(new_n737), .A4(new_n684), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n580), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n495), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT108), .B(G57gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1332gat));
  INV_X1    g598(.A(new_n796), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n803), .B(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n802), .B(new_n805), .ZN(G1333gat));
  NOR3_X1   g605(.A1(new_n796), .A2(new_n590), .A3(new_n577), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n549), .B(KEYINPUT111), .Z(new_n808));
  NAND2_X1  g607(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n590), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n542), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT112), .B(G78gat), .Z(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(G1335gat));
  NOR2_X1   g613(.A1(new_n611), .A2(new_n794), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n750), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n763), .B2(new_n764), .ZN(new_n818));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818), .B2(new_n495), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n580), .A2(new_n737), .A3(new_n815), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n580), .A2(KEYINPUT51), .A3(new_n737), .A4(new_n815), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n742), .A2(new_n635), .A3(new_n750), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(G1336gat));
  INV_X1    g627(.A(new_n634), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n818), .B2(new_n721), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n721), .A2(G92gat), .A3(new_n684), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n823), .B2(new_n825), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n822), .A2(KEYINPUT113), .A3(new_n824), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n836), .A3(new_n821), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n837), .A3(new_n831), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n830), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n839), .B2(new_n833), .ZN(G1337gat));
  OAI21_X1  g639(.A(G99gat), .B1(new_n818), .B2(new_n577), .ZN(new_n841));
  INV_X1    g640(.A(new_n549), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n842), .A2(G99gat), .A3(new_n684), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n826), .B2(new_n843), .ZN(G1338gat));
  OAI21_X1  g643(.A(G106gat), .B1(new_n818), .B2(new_n542), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n684), .A2(new_n542), .A3(G106gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n823), .B2(new_n825), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n835), .A2(new_n837), .A3(new_n846), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n845), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n848), .ZN(G1339gat));
  NOR2_X1   g651(.A1(new_n685), .A2(new_n794), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n697), .A2(new_n698), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n704), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n713), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n661), .A2(new_n858), .A3(new_n663), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n646), .A2(new_n595), .A3(new_n648), .ZN(new_n861));
  INV_X1    g660(.A(new_n670), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n672), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n649), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n675), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n682), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n675), .A3(new_n864), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n683), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT55), .B1(new_n867), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n867), .A2(new_n869), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT55), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n876), .A2(KEYINPUT114), .A3(new_n683), .A4(new_n870), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n859), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n749), .B1(new_n873), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n857), .A2(new_n684), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n664), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n611), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n853), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n464), .A3(new_n463), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n742), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n541), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT115), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(KEYINPUT115), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n749), .A2(G113gat), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT116), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n884), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n842), .A2(new_n495), .A3(new_n541), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n542), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G113gat), .B1(new_n895), .B2(new_n715), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(G1340gat));
  NAND2_X1  g696(.A1(new_n750), .A2(new_n212), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT117), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n888), .A2(new_n889), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G120gat), .B1(new_n895), .B2(new_n684), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1341gat));
  NAND2_X1  g701(.A1(new_n233), .A2(new_n234), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n895), .A2(new_n903), .A3(new_n738), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n611), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n903), .B2(new_n907), .ZN(G1342gat));
  NOR2_X1   g707(.A1(new_n664), .A2(new_n541), .ZN(new_n909));
  INV_X1    g708(.A(G134gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n886), .A2(KEYINPUT56), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G134gat), .B1(new_n895), .B2(new_n664), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT56), .B1(new_n886), .B2(new_n911), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G1343gat));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(new_n457), .C1(new_n853), .C2(new_n883), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n729), .A2(new_n495), .A3(new_n541), .ZN(new_n918));
  INV_X1    g717(.A(new_n853), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT119), .B1(new_n871), .B2(new_n872), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n876), .A2(new_n921), .A3(new_n683), .A4(new_n870), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n920), .A2(new_n710), .A3(new_n714), .A4(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n881), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n737), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n738), .B1(new_n925), .B2(new_n878), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n542), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n917), .B(new_n918), .C1(new_n927), .C2(new_n916), .ZN(new_n928));
  OAI21_X1  g727(.A(G141gat), .B1(new_n928), .B2(new_n715), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n884), .A2(new_n542), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n930), .A2(new_n391), .A3(new_n739), .A4(new_n918), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT120), .A4(new_n932), .ZN(new_n936));
  OAI21_X1  g735(.A(G141gat), .B1(new_n928), .B2(new_n749), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(new_n931), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n935), .B(new_n936), .C1(new_n932), .C2(new_n938), .ZN(G1344gat));
  NOR3_X1   g738(.A1(new_n859), .A2(new_n872), .A3(new_n871), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT121), .B1(new_n925), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n738), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n940), .A3(KEYINPUT121), .ZN(new_n943));
  OAI22_X1  g742(.A1(new_n942), .A2(new_n943), .B1(new_n739), .B2(new_n685), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n542), .A2(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT57), .B1(new_n884), .B2(new_n542), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n946), .A2(new_n750), .A3(new_n947), .A4(new_n918), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G148gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n389), .A2(KEYINPUT59), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n928), .B2(new_n684), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT122), .B1(new_n949), .B2(KEYINPUT59), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n918), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n750), .A2(new_n389), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n956), .ZN(G1345gat));
  OAI21_X1  g756(.A(new_n383), .B1(new_n955), .B2(new_n738), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n611), .A2(G155gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n928), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(G1346gat));
  NOR2_X1   g760(.A1(new_n928), .A2(new_n664), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n384), .B1(new_n962), .B2(KEYINPUT123), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(KEYINPUT123), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n729), .A2(new_n495), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n930), .A2(new_n384), .A3(new_n909), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1347gat));
  NOR2_X1   g766(.A1(new_n721), .A2(new_n742), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n893), .A2(new_n542), .A3(new_n808), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(G169gat), .B1(new_n969), .B2(new_n715), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n885), .A2(new_n968), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n794), .A2(new_n288), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT124), .ZN(G1348gat));
  NOR3_X1   g773(.A1(new_n969), .A2(new_n250), .A3(new_n684), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n885), .A2(new_n750), .A3(new_n968), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n250), .B2(new_n976), .ZN(G1349gat));
  OAI21_X1  g776(.A(G183gat), .B1(new_n969), .B2(new_n738), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n611), .A2(new_n265), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n971), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n969), .B2(new_n664), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n737), .A2(new_n264), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n984), .A2(new_n985), .B1(new_n971), .B2(new_n986), .ZN(G1351gat));
  AND2_X1   g786(.A1(new_n946), .A2(new_n947), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n577), .A2(new_n968), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n375), .B1(new_n991), .B2(new_n739), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n930), .A2(new_n989), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n993), .A2(G197gat), .A3(new_n749), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n992), .A2(new_n994), .ZN(G1352gat));
  NOR3_X1   g794(.A1(new_n993), .A2(G204gat), .A3(new_n684), .ZN(new_n996));
  XNOR2_X1  g795(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n996), .B(new_n997), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n988), .A2(new_n750), .A3(new_n990), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n376), .B2(new_n999), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n988), .A2(new_n611), .A3(new_n990), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(G211gat), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n611), .A2(new_n359), .ZN(new_n1004));
  OAI22_X1  g803(.A1(new_n1002), .A2(new_n1003), .B1(new_n993), .B2(new_n1004), .ZN(G1354gat));
  NAND3_X1  g804(.A1(new_n991), .A2(G218gat), .A3(new_n737), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n360), .B1(new_n993), .B2(new_n664), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1355gat));
endmodule


