//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(KEYINPUT98), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  AND2_X1   g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT9), .ZN(new_n210));
  XOR2_X1   g009(.A(G57gat), .B(G64gat), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G71gat), .B(G78gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(new_n217), .B(KEYINPUT102), .Z(new_n218));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G231gat), .ZN(new_n223));
  INV_X1    g022(.A(G233gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(G231gat), .A3(G233gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G155gat), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n228), .B(G211gat), .Z(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n217), .A2(new_n219), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n232), .B(new_n233), .Z(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n226), .B2(new_n227), .ZN(new_n236));
  OR3_X1    g035(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n231), .B2(new_n236), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT96), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OR3_X1    g041(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n241), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G29gat), .ZN(new_n246));
  INV_X1    g045(.A(G36gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G43gat), .B(G50gat), .Z(new_n249));
  INV_X1    g048(.A(KEYINPUT15), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT97), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n240), .B2(new_n243), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n249), .A2(new_n250), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT17), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G85gat), .A2(G92gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT7), .ZN(new_n263));
  INV_X1    g062(.A(G99gat), .ZN(new_n264));
  INV_X1    g063(.A(G106gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT8), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n263), .B(new_n266), .C1(G85gat), .C2(G92gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(G99gat), .B(G106gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT106), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G232gat), .A2(G233gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT103), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n257), .A2(new_n269), .B1(KEYINPUT41), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT106), .A3(new_n270), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n276), .A2(KEYINPUT41), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT107), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(G134gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G162gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n282), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n273), .A2(new_n288), .A3(new_n277), .A4(new_n278), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n283), .B2(new_n289), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G230gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(new_n224), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n269), .B(new_n217), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT10), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n218), .A2(new_n297), .A3(new_n270), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n296), .A2(new_n295), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G120gat), .B(G148gat), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G204gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n239), .A2(new_n292), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT35), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G113gat), .ZN(new_n318));
  INV_X1    g117(.A(G113gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G120gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT1), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G127gat), .A2(G134gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n326), .B(KEYINPUT69), .C1(new_n327), .C2(KEYINPUT1), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n320), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n320), .B2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n322), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT2), .ZN(new_n338));
  INV_X1    g137(.A(G148gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(G141gat), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(G148gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n344), .A2(KEYINPUT78), .A3(new_n337), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT78), .B1(new_n344), .B2(new_n337), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT79), .B1(new_n341), .B2(G148gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(new_n339), .A3(G141gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n341), .A2(G148gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT80), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n344), .A2(new_n356), .A3(new_n337), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n352), .A2(new_n338), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n336), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n329), .A2(new_n335), .A3(new_n347), .A4(new_n358), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n315), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT83), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n315), .ZN(new_n366));
  AND4_X1   g165(.A1(new_n329), .A2(new_n335), .A3(new_n347), .A4(new_n358), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n329), .A2(new_n335), .B1(new_n347), .B2(new_n358), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n363), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(new_n347), .B2(new_n358), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n336), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n347), .A2(new_n358), .A3(new_n373), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n374), .B2(new_n375), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n319), .A2(G120gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n317), .A2(G113gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(KEYINPUT70), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT1), .B1(new_n385), .B2(new_n332), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n386), .A2(new_n322), .B1(new_n323), .B2(new_n328), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n347), .A2(new_n358), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT4), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n380), .A2(new_n366), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT84), .B1(new_n372), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT81), .B1(new_n388), .B2(new_n373), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(new_n336), .A3(new_n376), .A4(new_n378), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(new_n315), .A3(new_n382), .A4(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n365), .A4(new_n371), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n315), .A3(new_n364), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT85), .B1(new_n382), .B2(new_n389), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n389), .A3(KEYINPUT85), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(G85gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n405), .A2(new_n410), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n403), .B1(new_n392), .B2(new_n397), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n415), .B2(new_n409), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n409), .B1(new_n398), .B2(new_n404), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G211gat), .B(G218gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT76), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  INV_X1    g222(.A(G197gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n306), .ZN(new_n425));
  NAND2_X1  g224(.A1(G197gat), .A2(G204gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT22), .ZN(new_n427));
  NAND2_X1  g226(.A1(G211gat), .A2(G218gat), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n425), .A2(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n429), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n422), .A2(KEYINPUT75), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G169gat), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n437), .A2(new_n304), .A3(KEYINPUT64), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT64), .B1(new_n437), .B2(new_n304), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT23), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(G169gat), .A2(G176gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT23), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT65), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT24), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT24), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(KEYINPUT65), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G190gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT66), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT66), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G190gat), .ZN(new_n455));
  AOI21_X1  g254(.A(G183gat), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n440), .B(new_n445), .C1(new_n451), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT25), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT26), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n438), .B2(new_n439), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n461), .A2(new_n441), .A3(KEYINPUT68), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT68), .B1(new_n461), .B2(new_n441), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n446), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n454), .A2(G190gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n452), .A2(KEYINPUT66), .ZN(new_n467));
  NOR2_X1   g266(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n468));
  AND2_X1   g267(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n466), .A2(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n465), .B1(new_n470), .B2(KEYINPUT28), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472));
  OR3_X1    g271(.A1(new_n472), .A2(new_n221), .A3(KEYINPUT27), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT28), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n455), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT27), .B1(new_n472), .B2(new_n221), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n464), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT25), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n465), .A2(new_n449), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n221), .A2(new_n452), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT24), .A3(new_n446), .ZN(new_n482));
  AND4_X1   g281(.A1(new_n479), .A2(new_n480), .A3(new_n482), .A4(new_n445), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n441), .A2(KEYINPUT23), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n458), .A2(new_n478), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n436), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n457), .A2(KEYINPUT25), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n435), .B1(new_n489), .B2(new_n478), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n434), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n436), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n489), .B2(new_n478), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n433), .C1(new_n493), .C2(new_n436), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G64gat), .B(G92gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT77), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G8gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(new_n247), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n495), .B2(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n499), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(new_n491), .A3(new_n502), .A4(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n420), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(G22gat), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n422), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n431), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n422), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n429), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n514), .B(new_n487), .C1(new_n516), .C2(new_n513), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n359), .B1(new_n518), .B2(KEYINPUT3), .ZN(new_n519));
  NAND2_X1  g318(.A1(G228gat), .A2(G233gat), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n378), .A2(new_n487), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT89), .B1(new_n433), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n433), .A2(new_n521), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n519), .A2(new_n520), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n433), .A2(new_n487), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n388), .B1(new_n527), .B2(new_n373), .ZN(new_n528));
  OAI211_X1 g327(.A(G228gat), .B(G233gat), .C1(new_n528), .C2(new_n523), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G50gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n526), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n511), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n526), .A2(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n530), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n510), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n486), .B2(new_n336), .ZN(new_n541));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n486), .A2(new_n336), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n489), .A2(KEYINPUT71), .A3(new_n387), .A4(new_n478), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT34), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n547));
  INV_X1    g346(.A(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT72), .B(G71gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G99gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G43gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n549), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT32), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT33), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n554), .B1(new_n549), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n546), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n553), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n545), .B(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n549), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n564), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT74), .A4(new_n569), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n572), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n539), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n314), .B1(new_n508), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n507), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT87), .B1(new_n418), .B2(KEYINPUT6), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n581));
  NOR4_X1   g380(.A1(new_n415), .A2(new_n412), .A3(new_n581), .A4(new_n409), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI211_X1 g382(.A(new_n410), .B(new_n403), .C1(new_n392), .C2(new_n397), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT86), .B1(new_n584), .B2(KEYINPUT6), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n398), .A2(new_n409), .A3(new_n404), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT86), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n581), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n414), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n579), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n564), .A2(new_n570), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n539), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(new_n314), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n491), .A2(new_n596), .A3(new_n494), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n491), .B2(new_n494), .ZN(new_n598));
  NOR4_X1   g397(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT38), .A4(new_n505), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n597), .A2(new_n598), .A3(new_n505), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n598), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n491), .A2(new_n596), .A3(new_n494), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n499), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT92), .A3(KEYINPUT38), .ZN(new_n607));
  AOI211_X1 g406(.A(new_n500), .B(new_n599), .C1(new_n603), .C2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n583), .A2(new_n608), .A3(new_n417), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n534), .A2(new_n538), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT91), .B(KEYINPUT39), .Z(new_n611));
  INV_X1    g410(.A(KEYINPUT85), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n390), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n394), .A3(new_n401), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(KEYINPUT90), .A3(new_n366), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT90), .B1(new_n614), .B2(new_n366), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n366), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n367), .A2(new_n368), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(new_n315), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n615), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n618), .A2(new_n625), .A3(KEYINPUT40), .A4(new_n409), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n626), .A2(new_n414), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n618), .A2(new_n625), .A3(new_n409), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n507), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n610), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n609), .A2(KEYINPUT93), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT93), .B1(new_n609), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n585), .A2(new_n414), .A3(new_n588), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n413), .A2(new_n419), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n507), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n572), .A2(new_n639), .A3(new_n574), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n637), .A2(new_n610), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n595), .B1(new_n634), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n208), .B1(new_n253), .B2(new_n256), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n261), .B2(new_n208), .ZN(new_n644));
  NAND2_X1  g443(.A1(G229gat), .A2(G233gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT18), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n257), .B(new_n208), .Z(new_n648));
  XOR2_X1   g447(.A(new_n645), .B(KEYINPUT13), .Z(new_n649));
  AOI22_X1  g448(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n651));
  INV_X1    g450(.A(new_n645), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n652), .B(new_n643), .C1(new_n261), .C2(new_n208), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n644), .A2(new_n651), .A3(KEYINPUT18), .A4(new_n645), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G169gat), .B(G197gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT18), .B1(new_n644), .B2(new_n645), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n665), .B2(KEYINPUT100), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n261), .A2(new_n208), .ZN(new_n668));
  INV_X1    g467(.A(new_n643), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n668), .A2(KEYINPUT18), .A3(new_n645), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n655), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n672), .B(new_n650), .C1(new_n674), .C2(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT101), .B1(new_n642), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n603), .A2(new_n607), .ZN(new_n680));
  INV_X1    g479(.A(new_n599), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n501), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n420), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n628), .A2(new_n629), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n684), .A2(new_n414), .A3(new_n579), .A4(new_n626), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n539), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n679), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n637), .A2(new_n610), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n640), .A2(new_n638), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n609), .A2(new_n631), .A3(KEYINPUT93), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n576), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n694), .A2(new_n539), .A3(new_n420), .A4(new_n507), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n695), .A2(new_n314), .B1(new_n590), .B2(new_n593), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n676), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n313), .B1(new_n678), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n583), .A2(new_n589), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  INV_X1    g503(.A(new_n313), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n698), .B1(new_n697), .B2(new_n676), .ZN(new_n706));
  AOI211_X1 g505(.A(KEYINPUT101), .B(new_n677), .C1(new_n691), .C2(new_n696), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n579), .B(new_n705), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT108), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n678), .A2(new_n699), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n579), .A4(new_n705), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT16), .B(G8gat), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n202), .A2(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n579), .A4(new_n714), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(KEYINPUT109), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1325gat));
  AOI21_X1  g523(.A(G15gat), .B1(new_n700), .B2(new_n694), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n640), .A2(new_n638), .A3(G15gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n700), .B2(new_n726), .ZN(G1326gat));
  NAND2_X1  g526(.A1(new_n700), .A2(new_n610), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT43), .B(G22gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  NAND2_X1  g529(.A1(new_n283), .A2(new_n289), .ZN(new_n731));
  INV_X1    g530(.A(new_n287), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n239), .A2(new_n311), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n710), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n246), .A3(new_n702), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n697), .A2(new_n735), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n697), .A2(new_n735), .B1(KEYINPUT110), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n676), .B(new_n736), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n701), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n747), .ZN(G1328gat));
  NOR3_X1   g547(.A1(new_n737), .A2(G36gat), .A3(new_n507), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G36gat), .B1(new_n746), .B2(new_n507), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1329gat));
  INV_X1    g552(.A(new_n694), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n737), .A2(G43gat), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G43gat), .B1(new_n746), .B2(new_n689), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1330gat));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n738), .A2(new_n761), .A3(new_n610), .ZN(new_n762));
  OAI21_X1  g561(.A(G50gat), .B1(new_n746), .B2(new_n539), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1331gat));
  NOR2_X1   g565(.A1(new_n642), .A2(new_n676), .ZN(new_n767));
  INV_X1    g566(.A(new_n239), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n768), .A2(new_n735), .A3(new_n312), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n702), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n507), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n776), .B(new_n777), .Z(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n770), .B2(new_n689), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n770), .A2(G71gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n754), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g581(.A1(new_n770), .A2(new_n539), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT113), .B(G78gat), .Z(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1335gat));
  NOR2_X1   g584(.A1(new_n239), .A2(new_n676), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT51), .B1(new_n741), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n697), .A2(new_n789), .A3(new_n735), .A4(new_n786), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n788), .A2(new_n311), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n702), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n311), .B(new_n786), .C1(new_n743), .C2(new_n745), .ZN(new_n793));
  INV_X1    g592(.A(G85gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n794), .A3(new_n701), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n792), .A2(new_n795), .ZN(G1336gat));
  NAND4_X1  g595(.A1(new_n788), .A2(new_n579), .A3(new_n311), .A4(new_n790), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n797), .A2(KEYINPUT115), .A3(G92gat), .ZN(new_n798));
  OAI21_X1  g597(.A(G92gat), .B1(new_n793), .B2(new_n507), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n797), .B2(G92gat), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n797), .A2(G92gat), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n803), .A2(KEYINPUT114), .A3(new_n799), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n803), .B2(KEYINPUT114), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n264), .A3(new_n694), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n793), .B2(new_n689), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n265), .A3(new_n610), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n793), .B2(new_n539), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n299), .B1(new_n297), .B2(new_n296), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n294), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n300), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n307), .B1(new_n300), .B2(KEYINPUT54), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n819), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n309), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n667), .B2(new_n675), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n672), .A2(new_n663), .A3(new_n650), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n644), .A2(new_n645), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n648), .A2(new_n649), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n662), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n825), .A2(new_n311), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n292), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n825), .A2(new_n828), .ZN(new_n831));
  INV_X1    g630(.A(new_n823), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n735), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n239), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n313), .A2(new_n676), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n577), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n702), .A3(new_n837), .A4(new_n507), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n677), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n702), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n840), .A2(new_n579), .A3(new_n592), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n319), .A3(new_n676), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(G1340gat));
  OAI21_X1  g642(.A(G120gat), .B1(new_n838), .B2(new_n312), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n317), .A3(new_n311), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n841), .B2(new_n239), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n838), .A2(new_n768), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g648(.A(G134gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n841), .A2(new_n850), .A3(new_n735), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n838), .B2(new_n292), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT116), .ZN(G1343gat));
  OAI21_X1  g655(.A(new_n610), .B1(new_n834), .B2(new_n835), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n610), .C1(new_n834), .C2(new_n835), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n702), .A2(new_n689), .A3(new_n507), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n676), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT118), .B(new_n702), .C1(new_n834), .C2(new_n835), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n689), .A2(new_n610), .A3(new_n507), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n870), .A2(new_n341), .A3(new_n676), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n865), .A2(new_n866), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT119), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n871), .B1(new_n868), .B2(new_n869), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n341), .A4(new_n676), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n861), .B2(new_n863), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT117), .B(new_n862), .C1(new_n859), .C2(new_n860), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n676), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n879), .B1(G141gat), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n874), .B1(new_n884), .B2(new_n866), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n876), .A2(new_n339), .A3(new_n311), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n311), .B1(new_n881), .B2(new_n882), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(G148gat), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n890));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n292), .B2(new_n823), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n735), .A2(KEYINPUT122), .A3(new_n832), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n831), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n830), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n835), .B1(new_n895), .B2(new_n768), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n858), .B1(new_n896), .B2(new_n539), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n899), .B(new_n858), .C1(new_n896), .C2(new_n539), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n860), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n862), .A2(KEYINPUT121), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n862), .A2(KEYINPUT121), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n901), .A2(new_n311), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n890), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n905), .ZN(G1345gat));
  INV_X1    g705(.A(new_n876), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n768), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n239), .B1(new_n881), .B2(new_n882), .ZN(new_n909));
  MUX2_X1   g708(.A(new_n908), .B(new_n909), .S(G155gat), .Z(G1346gat));
  OAI21_X1  g709(.A(new_n735), .B1(new_n881), .B2(new_n882), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n913), .B(new_n735), .C1(new_n881), .C2(new_n882), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(G162gat), .A3(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n292), .A2(G162gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n907), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n702), .A2(new_n507), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n836), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n591), .A3(new_n539), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n437), .A3(new_n676), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n837), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n677), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1348gat));
  NOR3_X1   g724(.A1(new_n923), .A2(new_n304), .A3(new_n312), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT125), .ZN(new_n927));
  AOI21_X1  g726(.A(G176gat), .B1(new_n921), .B2(new_n311), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n923), .B2(new_n768), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n919), .A2(KEYINPUT126), .A3(new_n837), .A4(new_n239), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(G183gat), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n921), .B(new_n239), .C1(new_n468), .C2(new_n469), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n923), .B2(new_n292), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n942), .B(G190gat), .C1(new_n923), .C2(new_n292), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n921), .A2(new_n475), .A3(new_n735), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(KEYINPUT127), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(G1351gat));
  INV_X1    g747(.A(new_n857), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n918), .A2(new_n689), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n949), .A2(new_n424), .A3(new_n676), .A4(new_n950), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n901), .A2(new_n676), .A3(new_n950), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n424), .ZN(G1352gat));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n954), .A2(G204gat), .A3(new_n312), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n901), .A2(new_n311), .A3(new_n950), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n306), .ZN(G1353gat));
  OR3_X1    g757(.A1(new_n954), .A2(G211gat), .A3(new_n768), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n901), .A2(new_n239), .A3(new_n950), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  NAND3_X1  g762(.A1(new_n901), .A2(new_n735), .A3(new_n950), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G218gat), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n292), .A2(G218gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n954), .B2(new_n966), .ZN(G1355gat));
endmodule


