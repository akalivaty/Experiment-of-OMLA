//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT66), .B(G2105), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n468), .B(G125), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(new_n473), .B2(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n464), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(KEYINPUT66), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(G137), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n469), .A2(new_n470), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n463), .A2(new_n473), .A3(KEYINPUT69), .A4(G137), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n475), .A2(new_n487), .ZN(G160));
  OAI221_X1 g063(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n464), .A2(new_n473), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n484), .B2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n473), .A2(KEYINPUT70), .A3(new_n476), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(G136), .B2(new_n496), .ZN(G162));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2104), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n469), .B2(new_n470), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n480), .A2(new_n482), .A3(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n505), .B2(new_n484), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n463), .A2(new_n473), .A3(new_n507), .A4(G138), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(G75), .A2(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(G651), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n518), .B2(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(G651), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n523), .A2(G50), .A3(G543), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n513), .A2(new_n514), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n523), .A2(G88), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(new_n525), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND2_X1  g104(.A1(new_n523), .A2(new_n524), .ZN(new_n530));
  INV_X1    g105(.A(new_n526), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n512), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n537), .A2(new_n538), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n521), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n532), .A2(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n534), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n532), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n534), .A2(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n521), .ZN(new_n553));
  AND3_X1   g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n531), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n532), .A2(G91), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  NAND3_X1  g142(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(G286));
  NAND4_X1  g143(.A1(new_n523), .A2(G87), .A3(new_n524), .A4(new_n526), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n519), .A2(new_n522), .B1(new_n518), .B2(G651), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n572), .A2(KEYINPUT73), .A3(G87), .A4(new_n526), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n523), .A2(G49), .A3(G543), .A4(new_n524), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G288));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n513), .B2(new_n514), .ZN(new_n580));
  AND2_X1   g155(.A1(G73), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n523), .A2(G48), .A3(G543), .A4(new_n524), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n523), .A2(G86), .A3(new_n524), .A4(new_n526), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n531), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n521), .B1(new_n588), .B2(KEYINPUT74), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(KEYINPUT74), .B2(new_n588), .ZN(new_n590));
  XNOR2_X1  g165(.A(KEYINPUT75), .B(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(G85), .A2(new_n532), .B1(new_n534), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(G290));
  NAND4_X1  g168(.A1(new_n523), .A2(G92), .A3(new_n524), .A4(new_n526), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n531), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n534), .A2(G54), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G171), .B2(new_n602), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(G171), .B2(new_n602), .ZN(G321));
  OR3_X1    g180(.A1(G168), .A2(KEYINPUT76), .A3(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT76), .B1(G168), .B2(new_n602), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n602), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(G297));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(G280));
  INV_X1    g185(.A(new_n601), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT77), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n616), .A2(KEYINPUT78), .B1(G868), .B2(new_n554), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(KEYINPUT78), .B2(new_n616), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n496), .A2(G135), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT80), .Z(new_n622));
  OR2_X1    g197(.A1(new_n463), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n484), .A2(new_n463), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n623), .A2(new_n625), .B1(new_n626), .B2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n473), .A2(new_n477), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n629), .A2(new_n630), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  NAND2_X1  g256(.A1(G160), .A2(G29), .ZN(new_n682));
  INV_X1    g257(.A(G34), .ZN(new_n683));
  AOI21_X1  g258(.A(G29), .B1(new_n683), .B2(KEYINPUT24), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(KEYINPUT24), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G2084), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G5), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G171), .B2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G1961), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n686), .A2(new_n687), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G32), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n496), .A2(G141), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n626), .A2(G129), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n702), .A2(new_n703), .B1(G105), .B2(new_n477), .ZN(new_n704));
  AND3_X1   g279(.A1(new_n698), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n697), .B1(new_n705), .B2(new_n696), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT27), .Z(new_n707));
  INV_X1    g282(.A(G1996), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n694), .B(new_n695), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G162), .A2(new_n696), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n696), .B2(G35), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2090), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n496), .A2(G139), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n719), .B(new_n722), .C1(new_n463), .C2(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G33), .B(new_n724), .S(G29), .Z(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(G2072), .Z(new_n726));
  INV_X1    g301(.A(G2090), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n715), .A2(new_n727), .A3(new_n716), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n696), .A2(G27), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n696), .ZN(new_n730));
  INV_X1    g305(.A(G2078), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n718), .A2(new_n726), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n711), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT30), .B(G28), .Z(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n689), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n689), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n738), .B1(new_n741), .B2(new_n742), .C1(new_n628), .C2(new_n696), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n691), .A2(G1961), .B1(new_n741), .B2(new_n742), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n696), .A2(KEYINPUT28), .A3(G26), .ZN(new_n749));
  AOI21_X1  g324(.A(KEYINPUT28), .B1(new_n696), .B2(G26), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n626), .A2(G128), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n496), .A2(G140), .ZN(new_n754));
  OAI221_X1 g329(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n749), .B(new_n750), .C1(new_n756), .C2(G29), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(G2067), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(G2067), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n689), .A2(G4), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n601), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1348), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n689), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n554), .B2(new_n689), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1341), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n760), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT87), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n689), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT23), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT90), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT89), .B(G1956), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n768), .B2(KEYINPUT87), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n734), .A2(new_n748), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n689), .A2(G23), .ZN(new_n778));
  INV_X1    g353(.A(G288), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n689), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n689), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n689), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n782), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n792));
  NOR2_X1   g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT83), .Z(new_n794));
  INV_X1    g369(.A(G119), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n792), .A2(new_n794), .B1(new_n491), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G131), .B2(new_n496), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT84), .Z(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n696), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n696), .A2(G25), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G24), .B(G290), .S(G16), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1986), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n802), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n791), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT85), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT85), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n810), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT36), .B1(new_n815), .B2(new_n808), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n777), .A2(new_n817), .ZN(G311));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n777), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n777), .B2(new_n817), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(G150));
  XOR2_X1   g397(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n572), .A2(G93), .A3(new_n526), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT93), .B(G55), .Z(new_n826));
  NAND3_X1  g401(.A1(new_n572), .A2(G543), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n827), .C1(new_n521), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n554), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(KEYINPUT94), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n828), .A2(new_n521), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(new_n834), .A3(new_n827), .A4(new_n825), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n830), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n837), .B1(new_n830), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n612), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n842), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n824), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n845), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n847), .A2(new_n823), .A3(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(G860), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT96), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT96), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n832), .A2(new_n835), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n724), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n756), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n496), .A2(G142), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n626), .A2(G130), .ZN(new_n863));
  OAI221_X1 g438(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n632), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n861), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n705), .B(G164), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n797), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n869), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(G160), .B(KEYINPUT97), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n628), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n875), .A3(new_n871), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g456(.A(G303), .B(G305), .Z(new_n882));
  XNOR2_X1  g457(.A(G290), .B(new_n779), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(KEYINPUT100), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G288), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n882), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT101), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT42), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n615), .A2(new_n840), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n615), .A2(new_n840), .ZN(new_n900));
  NAND2_X1  g475(.A1(G299), .A2(new_n601), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n561), .A2(new_n596), .A3(new_n565), .A4(new_n600), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT99), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n899), .B2(new_n900), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n905), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n905), .B2(new_n910), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n896), .A2(new_n898), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n896), .A2(new_n913), .A3(new_n898), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n855), .A2(new_n602), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n917), .ZN(G331));
  NAND2_X1  g494(.A1(new_n830), .A2(new_n836), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT95), .ZN(new_n921));
  OAI21_X1  g496(.A(G286), .B1(new_n545), .B2(new_n548), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n543), .B(KEYINPUT72), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n546), .A2(new_n547), .ZN(new_n924));
  NAND3_X1  g499(.A1(G168), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n830), .A2(new_n836), .A3(new_n837), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n921), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n925), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n838), .B2(new_n839), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n901), .A2(new_n933), .A3(new_n907), .A4(new_n902), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n906), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n931), .A2(KEYINPUT105), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT105), .B1(new_n931), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT103), .B1(new_n928), .B2(new_n930), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n840), .B2(new_n926), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n939), .A2(new_n941), .A3(new_n904), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n890), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n909), .B1(new_n939), .B2(new_n941), .ZN(new_n945));
  INV_X1    g520(.A(new_n903), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n928), .A2(new_n930), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n890), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n878), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n931), .A2(new_n935), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n931), .A2(KEYINPUT105), .A3(new_n935), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n893), .B1(new_n955), .B2(new_n942), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n878), .A4(new_n948), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n950), .A2(new_n958), .A3(KEYINPUT43), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n890), .B1(new_n945), .B2(new_n947), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT43), .B1(new_n949), .B2(new_n960), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n956), .A2(new_n878), .A3(new_n948), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n962), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  NAND3_X1  g545(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g548(.A1(G303), .A2(G8), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n977), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n972), .A2(new_n973), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT110), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n475), .A2(new_n487), .A3(G40), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n506), .A2(new_n508), .ZN(new_n984));
  INV_X1    g559(.A(new_n504), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G164), .B2(G1384), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n983), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n785), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n984), .B2(new_n985), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n983), .A3(new_n727), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n982), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n979), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n981), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n983), .A2(new_n993), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n574), .A2(G1976), .A3(new_n577), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(G8), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G305), .A2(G1981), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n583), .A2(new_n582), .A3(new_n584), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1009), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1012), .A2(new_n1004), .A3(G8), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n993), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n475), .A2(new_n487), .A3(G40), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1005), .B(G8), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT52), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1006), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1001), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1002), .A3(new_n779), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1009), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(G8), .A3(new_n1004), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n970), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n970), .C1(new_n1001), .C2(new_n1019), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n983), .A2(new_n988), .A3(new_n731), .A4(new_n990), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(KEYINPUT123), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT123), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n986), .B2(new_n987), .ZN(new_n1034));
  NOR3_X1   g609(.A1(G164), .A2(new_n989), .A3(G1384), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n1016), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(KEYINPUT53), .A4(new_n731), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n995), .A2(new_n983), .A3(new_n996), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n693), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT124), .B1(new_n1028), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(G171), .B1(new_n1033), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1032), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1030), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1028), .A2(new_n1041), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n693), .B2(new_n1039), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1048), .A3(G301), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1044), .A2(KEYINPUT54), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1016), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n993), .A2(KEYINPUT112), .A3(new_n994), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT112), .B1(new_n993), .B2(new_n994), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1051), .B(new_n727), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(new_n992), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT113), .B(new_n980), .C1(new_n1056), .C2(new_n982), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n982), .B1(new_n1055), .B2(new_n992), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n979), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n998), .A2(new_n1000), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1019), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1006), .A2(new_n1014), .A3(new_n1018), .A4(KEYINPUT114), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n981), .A2(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1050), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n991), .A2(new_n742), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n995), .A2(new_n983), .A3(new_n687), .A4(new_n996), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(KEYINPUT121), .A3(new_n1069), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(G168), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n982), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1070), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1074), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G286), .A2(G8), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(new_n1046), .A3(G301), .A4(new_n1042), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1067), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(G299), .B(KEYINPUT57), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1036), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n983), .A2(new_n996), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n995), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n1095), .B2(new_n1052), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1090), .B(new_n1092), .C1(new_n1096), .C2(G1956), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1098));
  INV_X1    g673(.A(G2067), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1039), .A2(new_n763), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n601), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1097), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1092), .B1(new_n1096), .B2(G1956), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1089), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT120), .B1(new_n1104), .B2(new_n1089), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1097), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1097), .A2(new_n1105), .A3(KEYINPUT61), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1100), .A2(new_n601), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1101), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT118), .B(G1996), .Z(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT58), .B(G1341), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n991), .A2(new_n1117), .B1(new_n1098), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n554), .ZN(new_n1120));
  NAND2_X1  g695(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1120), .A2(new_n1121), .B1(new_n1100), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1114), .A2(new_n1116), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1106), .B(new_n1108), .C1(new_n1113), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1027), .B1(new_n1088), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1068), .A2(KEYINPUT121), .A3(new_n1069), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT121), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1130), .A2(new_n1131), .A3(G286), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1076), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1081), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  AOI21_X1  g713(.A(G301), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1128), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1079), .A2(KEYINPUT62), .A3(new_n1081), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1061), .A2(new_n1066), .A3(new_n1139), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT125), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n980), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NOR4_X1   g724(.A1(new_n1077), .A2(new_n1019), .A3(new_n1149), .A4(G286), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1150), .A3(new_n1001), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1077), .A2(G286), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1061), .A2(new_n1066), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT115), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1061), .A2(new_n1066), .A3(KEYINPUT115), .A4(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1149), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1151), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1127), .A2(new_n1145), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n990), .A2(new_n1016), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n708), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT107), .ZN(new_n1162));
  INV_X1    g737(.A(new_n705), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n756), .B(new_n1099), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n708), .B2(new_n705), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1166), .B2(new_n1160), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n797), .B(new_n801), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1160), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(G290), .B(G1986), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1160), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1159), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(new_n798), .A3(new_n801), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(G2067), .B2(new_n756), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1176));
  NOR4_X1   g751(.A1(G290), .A2(G1986), .A3(new_n1016), .A4(new_n990), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1175), .A2(new_n1160), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1162), .B(KEYINPUT46), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n705), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1160), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT47), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1181), .A2(new_n1183), .A3(KEYINPUT47), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1186), .A2(KEYINPUT126), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1180), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT126), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1173), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g767(.A1(G401), .A2(G229), .A3(new_n461), .A4(G227), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n1194), .A3(new_n880), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


