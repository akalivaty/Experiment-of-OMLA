

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741;

  AND2_X2 U368 ( .A1(n738), .A2(KEYINPUT44), .ZN(n398) );
  XNOR2_X2 U369 ( .A(n376), .B(n375), .ZN(n552) );
  AND2_X2 U370 ( .A1(n543), .A2(n520), .ZN(n648) );
  XNOR2_X2 U371 ( .A(n479), .B(n478), .ZN(n517) );
  XNOR2_X2 U372 ( .A(n579), .B(n578), .ZN(n697) );
  AND2_X2 U373 ( .A1(n577), .A2(n576), .ZN(n579) );
  NOR2_X1 U374 ( .A1(n697), .A2(n580), .ZN(n581) );
  NOR2_X1 U375 ( .A1(n547), .A2(n549), .ZN(n531) );
  AND2_X1 U376 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U377 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U378 ( .A(n549), .B(KEYINPUT38), .ZN(n683) );
  XNOR2_X1 U379 ( .A(n510), .B(n509), .ZN(n666) );
  XNOR2_X1 U380 ( .A(n429), .B(n346), .ZN(n726) );
  INV_X2 U381 ( .A(G143), .ZN(n408) );
  OR2_X1 U382 ( .A1(n641), .A2(n655), .ZN(n575) );
  XNOR2_X1 U383 ( .A(n366), .B(KEYINPUT47), .ZN(n365) );
  NAND2_X1 U384 ( .A1(n349), .A2(n648), .ZN(n366) );
  XOR2_X1 U385 ( .A(KEYINPUT10), .B(n463), .Z(n495) );
  AND2_X1 U386 ( .A1(n344), .A2(KEYINPUT22), .ZN(n385) );
  NOR2_X1 U387 ( .A1(n666), .A2(n665), .ZN(n672) );
  INV_X1 U388 ( .A(KEYINPUT48), .ZN(n375) );
  XNOR2_X1 U389 ( .A(n495), .B(n368), .ZN(n367) );
  INV_X1 U390 ( .A(n494), .ZN(n368) );
  OR2_X1 U391 ( .A1(n536), .A2(n382), .ZN(n513) );
  XNOR2_X1 U392 ( .A(G469), .B(KEYINPUT69), .ZN(n488) );
  XNOR2_X1 U393 ( .A(n721), .B(n373), .ZN(n372) );
  INV_X1 U394 ( .A(KEYINPUT123), .ZN(n373) );
  XNOR2_X1 U395 ( .A(n405), .B(n404), .ZN(n403) );
  INV_X1 U396 ( .A(KEYINPUT86), .ZN(n404) );
  NAND2_X1 U397 ( .A1(n597), .A2(n596), .ZN(n405) );
  AND2_X1 U398 ( .A1(n396), .A2(n395), .ZN(n394) );
  AND2_X1 U399 ( .A1(n397), .A2(n585), .ZN(n389) );
  NAND2_X1 U400 ( .A1(n392), .A2(KEYINPUT85), .ZN(n391) );
  XNOR2_X1 U401 ( .A(n380), .B(KEYINPUT46), .ZN(n379) );
  AND2_X1 U402 ( .A1(n378), .A2(n377), .ZN(n355) );
  NOR2_X1 U403 ( .A1(n736), .A2(n741), .ZN(n380) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(G107), .Z(n431) );
  INV_X1 U405 ( .A(G146), .ZN(n452) );
  XNOR2_X1 U406 ( .A(n460), .B(n459), .ZN(n541) );
  XNOR2_X1 U407 ( .A(n458), .B(G475), .ZN(n459) );
  BUF_X1 U408 ( .A(n659), .Z(n720) );
  XNOR2_X1 U409 ( .A(G110), .B(G107), .ZN(n469) );
  INV_X1 U410 ( .A(KEYINPUT77), .ZN(n399) );
  NOR2_X1 U411 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U412 ( .A1(n683), .A2(n381), .ZN(n535) );
  NOR2_X1 U413 ( .A1(n570), .A2(n382), .ZN(n381) );
  BUF_X2 U414 ( .A(n517), .Z(n549) );
  XNOR2_X1 U415 ( .A(n519), .B(KEYINPUT19), .ZN(n369) );
  NAND2_X1 U416 ( .A1(n518), .A2(n682), .ZN(n519) );
  NAND2_X1 U417 ( .A1(n385), .A2(n383), .ZN(n384) );
  OR2_X1 U418 ( .A1(n344), .A2(KEYINPUT22), .ZN(n387) );
  BUF_X1 U419 ( .A(G953), .Z(n356) );
  XNOR2_X1 U420 ( .A(n505), .B(n367), .ZN(n711) );
  XNOR2_X1 U421 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U422 ( .A(n514), .B(n353), .ZN(n739) );
  INV_X1 U423 ( .A(KEYINPUT109), .ZN(n353) );
  AND2_X1 U424 ( .A1(n358), .A2(n357), .ZN(n641) );
  INV_X1 U425 ( .A(KEYINPUT101), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(G69) );
  XNOR2_X1 U427 ( .A(n725), .B(KEYINPUT124), .ZN(n370) );
  NAND2_X1 U428 ( .A1(n372), .A2(n724), .ZN(n371) );
  INV_X1 U429 ( .A(KEYINPUT60), .ZN(n362) );
  NOR2_X1 U430 ( .A1(n685), .A2(n665), .ZN(n344) );
  INV_X1 U431 ( .A(n534), .ZN(n382) );
  NOR2_X1 U432 ( .A1(n546), .A2(n640), .ZN(n345) );
  XOR2_X1 U433 ( .A(KEYINPUT4), .B(G131), .Z(n346) );
  NAND2_X1 U434 ( .A1(n454), .A2(n453), .ZN(n463) );
  AND2_X1 U435 ( .A1(n572), .A2(n534), .ZN(n347) );
  AND2_X1 U436 ( .A1(n401), .A2(n400), .ZN(n348) );
  BUF_X1 U437 ( .A(n569), .Z(n580) );
  NOR2_X1 U438 ( .A1(n687), .A2(n523), .ZN(n349) );
  INV_X1 U439 ( .A(n669), .ZN(n357) );
  NAND2_X1 U440 ( .A1(n608), .A2(n607), .ZN(n350) );
  XNOR2_X1 U441 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n351) );
  XOR2_X1 U442 ( .A(n610), .B(n609), .Z(n352) );
  INV_X1 U443 ( .A(KEYINPUT85), .ZN(n585) );
  XNOR2_X1 U444 ( .A(n613), .B(KEYINPUT91), .ZN(n714) );
  NOR2_X1 U445 ( .A1(n365), .A2(n739), .ZN(n524) );
  XNOR2_X2 U446 ( .A(n354), .B(n418), .ZN(n626) );
  XNOR2_X2 U447 ( .A(n487), .B(n413), .ZN(n354) );
  NAND2_X1 U448 ( .A1(n355), .A2(n379), .ZN(n376) );
  NAND2_X1 U449 ( .A1(n569), .A2(n563), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n531), .B(n351), .ZN(n532) );
  OR2_X2 U451 ( .A1(n541), .A2(n522), .ZN(n526) );
  XNOR2_X2 U452 ( .A(KEYINPUT94), .B(KEYINPUT17), .ZN(n464) );
  NAND2_X1 U453 ( .A1(n386), .A2(n384), .ZN(n595) );
  XNOR2_X1 U454 ( .A(n571), .B(n359), .ZN(n358) );
  NAND2_X1 U455 ( .A1(n575), .A2(n574), .ZN(n397) );
  XNOR2_X2 U456 ( .A(n360), .B(n399), .ZN(n664) );
  NAND2_X1 U457 ( .A1(n659), .A2(n601), .ZN(n360) );
  XNOR2_X1 U458 ( .A(n361), .B(n467), .ZN(n472) );
  XNOR2_X1 U459 ( .A(n466), .B(n468), .ZN(n361) );
  XNOR2_X1 U460 ( .A(n363), .B(n362), .ZN(G60) );
  NAND2_X1 U461 ( .A1(n638), .A2(n637), .ZN(n363) );
  XNOR2_X1 U462 ( .A(n364), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U463 ( .A1(n614), .A2(n637), .ZN(n364) );
  XNOR2_X1 U464 ( .A(n367), .B(n726), .ZN(n731) );
  AND2_X1 U465 ( .A1(n369), .A2(n374), .ZN(n520) );
  NAND2_X1 U466 ( .A1(n369), .A2(n559), .ZN(n562) );
  NAND2_X1 U467 ( .A1(n672), .A2(n374), .ZN(n570) );
  XNOR2_X2 U468 ( .A(n374), .B(KEYINPUT1), .ZN(n671) );
  NAND2_X1 U469 ( .A1(n543), .A2(n374), .ZN(n544) );
  XNOR2_X2 U470 ( .A(n489), .B(n488), .ZN(n374) );
  XNOR2_X1 U471 ( .A(n657), .B(n533), .ZN(n377) );
  XNOR2_X1 U472 ( .A(n524), .B(KEYINPUT74), .ZN(n378) );
  INV_X1 U473 ( .A(n569), .ZN(n383) );
  NAND2_X1 U474 ( .A1(n595), .A2(n564), .ZN(n586) );
  NAND2_X1 U475 ( .A1(n390), .A2(n389), .ZN(n396) );
  NOR2_X1 U476 ( .A1(n616), .A2(n398), .ZN(n390) );
  NOR2_X2 U477 ( .A1(n568), .A2(n666), .ZN(n616) );
  NAND2_X1 U478 ( .A1(n394), .A2(n391), .ZN(n599) );
  NAND2_X1 U479 ( .A1(n393), .A2(n397), .ZN(n392) );
  INV_X1 U480 ( .A(n616), .ZN(n393) );
  NAND2_X1 U481 ( .A1(n398), .A2(KEYINPUT85), .ZN(n395) );
  AND2_X4 U482 ( .A1(n664), .A2(n350), .ZN(n706) );
  INV_X4 U483 ( .A(G953), .ZN(n728) );
  NAND2_X1 U484 ( .A1(n403), .A2(n598), .ZN(n400) );
  NAND2_X1 U485 ( .A1(n402), .A2(KEYINPUT44), .ZN(n401) );
  INV_X1 U486 ( .A(n403), .ZN(n402) );
  BUF_X1 U487 ( .A(n706), .Z(n710) );
  XOR2_X1 U488 ( .A(n633), .B(n635), .Z(n406) );
  AND2_X1 U489 ( .A1(n450), .A2(G210), .ZN(n407) );
  INV_X1 U490 ( .A(KEYINPUT82), .ZN(n533) );
  INV_X1 U491 ( .A(KEYINPUT12), .ZN(n444) );
  XNOR2_X1 U492 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U493 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U494 ( .A(G134), .ZN(n409) );
  XNOR2_X1 U495 ( .A(n412), .B(n407), .ZN(n413) );
  INV_X1 U496 ( .A(KEYINPUT71), .ZN(n499) );
  XNOR2_X1 U497 ( .A(n500), .B(n499), .ZN(n501) );
  BUF_X1 U498 ( .A(n572), .Z(n669) );
  INV_X1 U499 ( .A(n714), .ZN(n637) );
  XNOR2_X2 U500 ( .A(n408), .B(G128), .ZN(n468) );
  XNOR2_X2 U501 ( .A(n468), .B(n409), .ZN(n429) );
  XNOR2_X2 U502 ( .A(n726), .B(G146), .ZN(n487) );
  XOR2_X1 U503 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n411) );
  XNOR2_X1 U504 ( .A(G137), .B(KEYINPUT75), .ZN(n410) );
  XNOR2_X1 U505 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U506 ( .A1(n356), .A2(G237), .ZN(n450) );
  XNOR2_X1 U507 ( .A(G119), .B(G116), .ZN(n415) );
  XNOR2_X1 U508 ( .A(G113), .B(KEYINPUT70), .ZN(n414) );
  XNOR2_X1 U509 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U510 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n416) );
  XNOR2_X1 U511 ( .A(n417), .B(n416), .ZN(n715) );
  XNOR2_X1 U512 ( .A(KEYINPUT67), .B(G101), .ZN(n482) );
  XNOR2_X1 U513 ( .A(n715), .B(n482), .ZN(n473) );
  INV_X1 U514 ( .A(n473), .ZN(n418) );
  INV_X1 U515 ( .A(G902), .ZN(n421) );
  NAND2_X1 U516 ( .A1(n626), .A2(n421), .ZN(n419) );
  XNOR2_X2 U517 ( .A(n419), .B(G472), .ZN(n572) );
  INV_X1 U518 ( .A(G237), .ZN(n420) );
  NAND2_X1 U519 ( .A1(n421), .A2(n420), .ZN(n476) );
  NAND2_X1 U520 ( .A1(n476), .A2(G214), .ZN(n682) );
  NAND2_X1 U521 ( .A1(n572), .A2(n682), .ZN(n422) );
  XNOR2_X1 U522 ( .A(n422), .B(KEYINPUT30), .ZN(n536) );
  NAND2_X1 U523 ( .A1(G234), .A2(G237), .ZN(n423) );
  XNOR2_X1 U524 ( .A(KEYINPUT14), .B(n423), .ZN(n425) );
  NAND2_X1 U525 ( .A1(G902), .A2(n425), .ZN(n554) );
  NOR2_X1 U526 ( .A1(G900), .A2(n554), .ZN(n424) );
  NAND2_X1 U527 ( .A1(n424), .A2(n356), .ZN(n427) );
  NAND2_X1 U528 ( .A1(G952), .A2(n425), .ZN(n695) );
  NOR2_X1 U529 ( .A1(n695), .A2(n356), .ZN(n426) );
  XNOR2_X1 U530 ( .A(n426), .B(KEYINPUT95), .ZN(n558) );
  NAND2_X1 U531 ( .A1(n427), .A2(n558), .ZN(n428) );
  XOR2_X1 U532 ( .A(n428), .B(KEYINPUT79), .Z(n534) );
  XNOR2_X1 U533 ( .A(KEYINPUT106), .B(KEYINPUT7), .ZN(n438) );
  INV_X1 U534 ( .A(n429), .ZN(n433) );
  XNOR2_X1 U535 ( .A(G116), .B(G122), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U537 ( .A(n433), .B(n432), .ZN(n436) );
  NAND2_X1 U538 ( .A1(G234), .A2(n728), .ZN(n434) );
  XOR2_X1 U539 ( .A(KEYINPUT8), .B(n434), .Z(n496) );
  NAND2_X1 U540 ( .A1(G217), .A2(n496), .ZN(n435) );
  XNOR2_X1 U541 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U542 ( .A(n438), .B(n437), .ZN(n707) );
  NOR2_X2 U543 ( .A1(n707), .A2(G902), .ZN(n439) );
  XNOR2_X2 U544 ( .A(n439), .B(G478), .ZN(n540) );
  XOR2_X1 U545 ( .A(G140), .B(KEYINPUT11), .Z(n441) );
  XNOR2_X1 U546 ( .A(G143), .B(G122), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n441), .B(n440), .ZN(n449) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n443) );
  XNOR2_X1 U549 ( .A(G131), .B(KEYINPUT102), .ZN(n442) );
  XNOR2_X1 U550 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U551 ( .A(G113), .B(G104), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n449), .B(n448), .ZN(n457) );
  NAND2_X1 U553 ( .A1(G214), .A2(n450), .ZN(n455) );
  INV_X1 U554 ( .A(G125), .ZN(n451) );
  NAND2_X1 U555 ( .A1(G146), .A2(n451), .ZN(n454) );
  NAND2_X1 U556 ( .A1(n452), .A2(G125), .ZN(n453) );
  XOR2_X1 U557 ( .A(n455), .B(n495), .Z(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n633) );
  NOR2_X1 U559 ( .A1(G902), .A2(n633), .ZN(n460) );
  XNOR2_X1 U560 ( .A(KEYINPUT13), .B(KEYINPUT105), .ZN(n458) );
  NOR2_X1 U561 ( .A1(n540), .A2(n541), .ZN(n461) );
  XNOR2_X1 U562 ( .A(n461), .B(KEYINPUT108), .ZN(n582) );
  XNOR2_X1 U563 ( .A(KEYINPUT18), .B(KEYINPUT4), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n467) );
  NAND2_X1 U565 ( .A1(n728), .A2(G224), .ZN(n465) );
  XNOR2_X1 U566 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n469), .B(G104), .ZN(n484) );
  XNOR2_X1 U568 ( .A(KEYINPUT16), .B(G122), .ZN(n470) );
  XNOR2_X1 U569 ( .A(n470), .B(KEYINPUT73), .ZN(n471) );
  XNOR2_X1 U570 ( .A(n484), .B(n471), .ZN(n716) );
  XNOR2_X1 U571 ( .A(n472), .B(n716), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n474), .B(n473), .ZN(n618) );
  XNOR2_X1 U573 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n475) );
  XNOR2_X1 U574 ( .A(n475), .B(G902), .ZN(n603) );
  NAND2_X1 U575 ( .A1(n618), .A2(n603), .ZN(n479) );
  NAND2_X1 U576 ( .A1(n476), .A2(G210), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n477), .B(KEYINPUT78), .ZN(n478) );
  INV_X1 U578 ( .A(n549), .ZN(n480) );
  NAND2_X1 U579 ( .A1(n582), .A2(n480), .ZN(n511) );
  NAND2_X1 U580 ( .A1(G227), .A2(n728), .ZN(n481) );
  XNOR2_X1 U581 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U582 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U583 ( .A(G137), .B(G140), .Z(n494) );
  XNOR2_X1 U584 ( .A(n485), .B(n494), .ZN(n486) );
  XNOR2_X1 U585 ( .A(n487), .B(n486), .ZN(n610) );
  NOR2_X1 U586 ( .A1(n610), .A2(G902), .ZN(n489) );
  NAND2_X1 U587 ( .A1(n603), .A2(G234), .ZN(n490) );
  XNOR2_X1 U588 ( .A(KEYINPUT20), .B(n490), .ZN(n506) );
  NAND2_X1 U589 ( .A1(G221), .A2(n506), .ZN(n493) );
  XOR2_X1 U590 ( .A(KEYINPUT100), .B(KEYINPUT21), .Z(n491) );
  XNOR2_X1 U591 ( .A(n491), .B(KEYINPUT99), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n493), .B(n492), .ZN(n665) );
  NAND2_X1 U593 ( .A1(n496), .A2(G221), .ZN(n504) );
  XOR2_X1 U594 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n498) );
  XNOR2_X1 U595 ( .A(G128), .B(KEYINPUT23), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n498), .B(n497), .ZN(n502) );
  XNOR2_X1 U597 ( .A(G119), .B(G110), .ZN(n500) );
  XNOR2_X1 U598 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U599 ( .A1(n711), .A2(G902), .ZN(n510) );
  NAND2_X1 U600 ( .A1(n506), .A2(G217), .ZN(n508) );
  XOR2_X1 U601 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n507) );
  XNOR2_X1 U602 ( .A(n508), .B(n507), .ZN(n509) );
  OR2_X1 U603 ( .A1(n511), .A2(n570), .ZN(n512) );
  NOR2_X1 U604 ( .A1(n513), .A2(n512), .ZN(n514) );
  INV_X1 U605 ( .A(n666), .ZN(n592) );
  NOR2_X1 U606 ( .A1(n592), .A2(n665), .ZN(n527) );
  NAND2_X1 U607 ( .A1(n527), .A2(n347), .ZN(n516) );
  INV_X1 U608 ( .A(KEYINPUT28), .ZN(n515) );
  XNOR2_X1 U609 ( .A(n516), .B(n515), .ZN(n543) );
  INV_X1 U610 ( .A(n517), .ZN(n518) );
  INV_X1 U611 ( .A(n540), .ZN(n522) );
  NAND2_X1 U612 ( .A1(n541), .A2(n522), .ZN(n521) );
  XOR2_X1 U613 ( .A(n521), .B(KEYINPUT107), .Z(n640) );
  NAND2_X1 U614 ( .A1(n640), .A2(n526), .ZN(n574) );
  INV_X1 U615 ( .A(n574), .ZN(n687) );
  INV_X1 U616 ( .A(KEYINPUT68), .ZN(n523) );
  INV_X1 U617 ( .A(n671), .ZN(n565) );
  INV_X1 U618 ( .A(KEYINPUT6), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n572), .B(n525), .ZN(n576) );
  NAND2_X1 U620 ( .A1(n682), .A2(n534), .ZN(n529) );
  INV_X2 U621 ( .A(n526), .ZN(n652) );
  NAND2_X1 U622 ( .A1(n652), .A2(n527), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n576), .A2(n530), .ZN(n547) );
  NOR2_X1 U624 ( .A1(n565), .A2(n532), .ZN(n657) );
  XNOR2_X1 U625 ( .A(n537), .B(KEYINPUT39), .ZN(n546) );
  NOR2_X1 U626 ( .A1(n546), .A2(n526), .ZN(n539) );
  XNOR2_X1 U627 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n538) );
  XNOR2_X1 U628 ( .A(n539), .B(n538), .ZN(n736) );
  NAND2_X1 U629 ( .A1(n683), .A2(n682), .ZN(n686) );
  NAND2_X1 U630 ( .A1(n541), .A2(n540), .ZN(n685) );
  NOR2_X1 U631 ( .A1(n686), .A2(n685), .ZN(n542) );
  XNOR2_X1 U632 ( .A(n542), .B(KEYINPUT41), .ZN(n696) );
  NOR2_X1 U633 ( .A1(n696), .A2(n544), .ZN(n545) );
  XNOR2_X1 U634 ( .A(n545), .B(KEYINPUT42), .ZN(n741) );
  OR2_X1 U635 ( .A1(n671), .A2(n547), .ZN(n548) );
  XNOR2_X1 U636 ( .A(KEYINPUT43), .B(n548), .ZN(n550) );
  AND2_X1 U637 ( .A1(n550), .A2(n549), .ZN(n615) );
  NOR2_X1 U638 ( .A1(n345), .A2(n615), .ZN(n551) );
  AND2_X2 U639 ( .A1(n552), .A2(n551), .ZN(n602) );
  NAND2_X1 U640 ( .A1(n602), .A2(KEYINPUT2), .ZN(n553) );
  XNOR2_X1 U641 ( .A(n553), .B(KEYINPUT81), .ZN(n601) );
  INV_X1 U642 ( .A(n554), .ZN(n555) );
  NOR2_X1 U643 ( .A1(G898), .A2(n728), .ZN(n718) );
  NAND2_X1 U644 ( .A1(n555), .A2(n718), .ZN(n556) );
  XNOR2_X1 U645 ( .A(n556), .B(KEYINPUT96), .ZN(n557) );
  NAND2_X1 U646 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U647 ( .A(KEYINPUT90), .B(KEYINPUT0), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n560), .B(KEYINPUT66), .ZN(n561) );
  XNOR2_X2 U649 ( .A(n562), .B(n561), .ZN(n569) );
  INV_X1 U650 ( .A(KEYINPUT22), .ZN(n563) );
  INV_X1 U651 ( .A(n576), .ZN(n564) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT83), .ZN(n566) );
  NAND2_X1 U653 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U654 ( .A(n567), .B(KEYINPUT84), .ZN(n568) );
  NOR2_X1 U655 ( .A1(n580), .A2(n570), .ZN(n571) );
  AND2_X1 U656 ( .A1(n672), .A2(n671), .ZN(n577) );
  AND2_X1 U657 ( .A1(n669), .A2(n577), .ZN(n678) );
  NAND2_X1 U658 ( .A1(n383), .A2(n678), .ZN(n573) );
  XNOR2_X1 U659 ( .A(n573), .B(KEYINPUT31), .ZN(n655) );
  XNOR2_X1 U660 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n578) );
  XNOR2_X1 U661 ( .A(n581), .B(KEYINPUT34), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X2 U663 ( .A(n584), .B(KEYINPUT35), .ZN(n738) );
  NOR2_X1 U664 ( .A1(n738), .A2(KEYINPUT44), .ZN(n598) );
  INV_X1 U665 ( .A(n586), .ZN(n588) );
  AND2_X1 U666 ( .A1(n671), .A2(n666), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n591) );
  INV_X1 U668 ( .A(KEYINPUT64), .ZN(n589) );
  XNOR2_X1 U669 ( .A(n589), .B(KEYINPUT32), .ZN(n590) );
  XNOR2_X1 U670 ( .A(n591), .B(n590), .ZN(n617) );
  INV_X1 U671 ( .A(n617), .ZN(n597) );
  OR2_X1 U672 ( .A1(n669), .A2(n592), .ZN(n593) );
  NOR2_X1 U673 ( .A1(n671), .A2(n593), .ZN(n594) );
  AND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n646) );
  INV_X1 U675 ( .A(n646), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n599), .A2(n348), .ZN(n600) );
  XNOR2_X2 U677 ( .A(n600), .B(KEYINPUT45), .ZN(n659) );
  INV_X1 U678 ( .A(n603), .ZN(n605) );
  AND2_X1 U679 ( .A1(n602), .A2(n605), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n659), .A2(n604), .ZN(n608) );
  INV_X1 U681 ( .A(KEYINPUT2), .ZN(n606) );
  OR2_X1 U682 ( .A1(n603), .A2(n606), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n706), .A2(G469), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n609) );
  XNOR2_X1 U685 ( .A(n611), .B(n352), .ZN(n614) );
  INV_X1 U686 ( .A(G952), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n612), .A2(n356), .ZN(n613) );
  XOR2_X1 U688 ( .A(n615), .B(G140), .Z(G42) );
  XOR2_X1 U689 ( .A(n616), .B(G101), .Z(G3) );
  XOR2_X1 U690 ( .A(n617), .B(G119), .Z(G21) );
  NAND2_X1 U691 ( .A1(n706), .A2(G210), .ZN(n622) );
  XNOR2_X1 U692 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n619) );
  XOR2_X1 U693 ( .A(n619), .B(KEYINPUT55), .Z(n620) );
  XNOR2_X1 U694 ( .A(n618), .B(n620), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U696 ( .A1(n623), .A2(n714), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n624), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U698 ( .A1(n706), .A2(G472), .ZN(n628) );
  XNOR2_X1 U699 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X2 U702 ( .A1(n629), .A2(n714), .ZN(n632) );
  XNOR2_X1 U703 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n630) );
  XOR2_X1 U704 ( .A(n630), .B(KEYINPUT88), .Z(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(G57) );
  NAND2_X1 U706 ( .A1(n706), .A2(G475), .ZN(n636) );
  XNOR2_X1 U707 ( .A(KEYINPUT65), .B(KEYINPUT122), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT59), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n636), .B(n406), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n641), .A2(n652), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n639), .B(G104), .ZN(G6) );
  XOR2_X1 U712 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n643) );
  INV_X1 U713 ( .A(n640), .ZN(n654) );
  NAND2_X1 U714 ( .A1(n641), .A2(n654), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n645) );
  XOR2_X1 U716 ( .A(G107), .B(KEYINPUT27), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U718 ( .A(G110), .B(n646), .Z(n647) );
  XNOR2_X1 U719 ( .A(KEYINPUT114), .B(n647), .ZN(G12) );
  XOR2_X1 U720 ( .A(G128), .B(KEYINPUT29), .Z(n650) );
  NAND2_X1 U721 ( .A1(n648), .A2(n654), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(G30) );
  NAND2_X1 U723 ( .A1(n648), .A2(n652), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n651), .B(G146), .ZN(G48) );
  NAND2_X1 U725 ( .A1(n655), .A2(n652), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(G113), .ZN(G15) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n656), .B(G116), .ZN(G18) );
  XNOR2_X1 U729 ( .A(G125), .B(n657), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U731 ( .A(G134), .B(n345), .Z(G36) );
  XOR2_X1 U732 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n705) );
  NOR2_X1 U733 ( .A1(n720), .A2(KEYINPUT2), .ZN(n662) );
  NOR2_X1 U734 ( .A1(n602), .A2(KEYINPUT2), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(KEYINPUT80), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n701) );
  XOR2_X1 U738 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n668) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n670), .A2(n357), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT50), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U745 ( .A(KEYINPUT117), .B(n676), .Z(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U747 ( .A(KEYINPUT51), .B(n679), .Z(n680) );
  NOR2_X1 U748 ( .A1(n696), .A2(n680), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(KEYINPUT118), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n697), .A2(n690), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U756 ( .A(n693), .B(KEYINPUT52), .ZN(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U761 ( .A(KEYINPUT119), .B(n702), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n703), .A2(n728), .ZN(n704) );
  XNOR2_X1 U763 ( .A(n705), .B(n704), .ZN(G75) );
  NAND2_X1 U764 ( .A1(n710), .A2(G478), .ZN(n708) );
  XNOR2_X1 U765 ( .A(n707), .B(n708), .ZN(n709) );
  NOR2_X1 U766 ( .A1(n714), .A2(n709), .ZN(G63) );
  NAND2_X1 U767 ( .A1(n710), .A2(G217), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U770 ( .A(n715), .B(G101), .ZN(n717) );
  XNOR2_X1 U771 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n720), .A2(n728), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n356), .A2(G224), .ZN(n722) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n722), .ZN(n723) );
  NAND2_X1 U776 ( .A1(n723), .A2(G898), .ZN(n724) );
  XNOR2_X1 U777 ( .A(n731), .B(n602), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n727), .B(KEYINPUT125), .ZN(n729) );
  NAND2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U780 ( .A(n730), .B(KEYINPUT126), .ZN(n735) );
  XNOR2_X1 U781 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U782 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U783 ( .A1(n733), .A2(n356), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n735), .A2(n734), .ZN(G72) );
  XNOR2_X1 U785 ( .A(G131), .B(n736), .ZN(n737) );
  XNOR2_X1 U786 ( .A(n737), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U787 ( .A(n738), .B(G122), .Z(G24) );
  XNOR2_X1 U788 ( .A(n739), .B(G143), .ZN(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(KEYINPUT115), .ZN(G45) );
  XOR2_X1 U790 ( .A(G137), .B(n741), .Z(G39) );
endmodule

