//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n598, new_n601, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1109, new_n1110;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n465), .A2(G112), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(new_n465), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n479), .B2(G124), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT69), .Z(G162));
  OAI211_X1 g056(.A(G138), .B(new_n465), .C1(new_n461), .C2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(new_n465), .A3(G138), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n463), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT71), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n483), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n478), .A2(G126), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n507));
  XOR2_X1   g082(.A(KEYINPUT6), .B(G651), .Z(new_n508));
  OAI22_X1  g083(.A1(new_n506), .A2(KEYINPUT72), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  NAND2_X1  g087(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(G543), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT74), .B(G51), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n503), .A2(new_n514), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n519), .A2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n523), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n529), .A2(new_n530), .B1(new_n517), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n505), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  INV_X1    g114(.A(new_n523), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT77), .B(G81), .Z(new_n541));
  AOI22_X1  g116(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n513), .A2(G543), .A3(new_n516), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G43), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT76), .B1(new_n537), .B2(new_n505), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT80), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n543), .A2(G53), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT81), .A2(KEYINPUT9), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n505), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n523), .B(KEYINPUT82), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  NAND2_X1  g140(.A1(new_n562), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n543), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n562), .A2(G86), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n503), .A2(G61), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n505), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n570), .A2(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n543), .A2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n505), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n540), .A2(G85), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n562), .A2(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(new_n503), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n543), .A2(G54), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n583), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n583), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT83), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(G868), .B2(new_n598), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(G868), .B2(new_n598), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G860), .ZN(G148));
  OAI21_X1  g177(.A(G868), .B1(new_n592), .B2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n464), .A2(G135), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n465), .A2(G111), .ZN(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n479), .B2(G123), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT84), .Z(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND2_X1  g187(.A1(new_n488), .A2(new_n466), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT13), .B(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(KEYINPUT14), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT87), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT86), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2451), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n626), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n633), .A2(G14), .A3(new_n634), .ZN(G401));
  XNOR2_X1  g210(.A(G2084), .B(G2090), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT88), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(G2072), .A2(G2078), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n442), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT17), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n638), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT90), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n640), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n637), .B(new_n646), .C1(new_n641), .C2(new_n643), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT89), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n637), .A2(new_n643), .A3(new_n640), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2096), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT20), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n656), .B2(new_n660), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n656), .A2(KEYINPUT92), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  MUX2_X1   g248(.A(G6), .B(G305), .S(G16), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT32), .B(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(G166), .A2(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G16), .B2(G22), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n683), .B2(G23), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT33), .B(G1976), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n680), .B(new_n681), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n676), .B(new_n687), .C1(new_n685), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n683), .A2(G24), .ZN(new_n692));
  INV_X1    g267(.A(G290), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n683), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G1986), .Z(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  INV_X1    g273(.A(G107), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G2105), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G131), .B2(new_n464), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n479), .A2(G119), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n697), .B1(new_n705), .B2(new_n696), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n690), .A2(new_n691), .A3(new_n695), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT36), .ZN(new_n710));
  NOR2_X1   g285(.A1(G29), .A2(G33), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT95), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n488), .A2(G127), .ZN(new_n715));
  NAND2_X1  g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n465), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n714), .B(new_n717), .C1(G139), .C2(new_n464), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT96), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n712), .B1(new_n720), .B2(new_n696), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2072), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n724), .B2(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(KEYINPUT24), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n472), .B2(new_n696), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n479), .A2(G129), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT26), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n731), .A2(new_n732), .B1(G105), .B2(new_n466), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n464), .A2(G141), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT97), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G29), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(G29), .B2(G32), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n741), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT99), .Z(new_n747));
  OAI221_X1 g322(.A(new_n722), .B1(new_n723), .B2(new_n727), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n696), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n696), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT104), .ZN(new_n754));
  NOR2_X1   g329(.A1(G168), .A2(new_n683), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n683), .B2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT102), .B(KEYINPUT31), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G11), .Z(new_n760));
  AND2_X1   g335(.A1(new_n727), .A2(new_n723), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT103), .B(G28), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT30), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(KEYINPUT30), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n760), .B(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n758), .B(new_n765), .C1(new_n696), .C2(new_n611), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n745), .B2(new_n747), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n756), .A2(new_n757), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT101), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n683), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n683), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1961), .Z(new_n772));
  AND4_X1   g347(.A1(new_n754), .A2(new_n767), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n750), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n749), .B2(new_n748), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT105), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n696), .A2(G35), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT106), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n696), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT29), .B(G2090), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n683), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n547), .B2(new_n683), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n696), .A2(G26), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n479), .A2(G128), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n464), .A2(G140), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n465), .A2(G116), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n788), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2067), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n783), .A2(new_n786), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n683), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n593), .B2(new_n683), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1348), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n683), .A2(G20), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT23), .Z(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n796), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n710), .A2(new_n777), .A3(new_n778), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NOR2_X1   g382(.A1(new_n592), .A2(new_n601), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  INV_X1    g384(.A(G67), .ZN(new_n810));
  INV_X1    g385(.A(G80), .ZN(new_n811));
  INV_X1    g386(.A(G543), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n588), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT107), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT107), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n815), .B1(new_n811), .B2(new_n812), .C1(new_n588), .C2(new_n810), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n814), .A2(G651), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n543), .A2(G55), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n540), .A2(G93), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n547), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n546), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n809), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  INV_X1    g401(.A(G860), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n822), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n720), .B(new_n737), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n704), .B(new_n614), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT108), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n484), .B1(new_n463), .B2(new_n486), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n490), .ZN(new_n838));
  AOI221_X4 g413(.A(new_n836), .B1(new_n482), .B2(KEYINPUT4), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT108), .B1(new_n840), .B2(new_n483), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n500), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n793), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n464), .A2(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n465), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n479), .B2(G130), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n835), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n611), .B(new_n472), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT109), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n854), .B(new_n855), .C1(new_n852), .C2(new_n850), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g432(.A(G303), .B(G305), .ZN(new_n858));
  XNOR2_X1  g433(.A(G288), .B(G290), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT42), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n598), .B(new_n592), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n592), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n824), .ZN(new_n866));
  MUX2_X1   g441(.A(new_n862), .B(new_n864), .S(new_n866), .Z(new_n867));
  AOI21_X1  g442(.A(new_n861), .B1(new_n867), .B2(KEYINPUT110), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT110), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(G868), .B2(new_n820), .ZN(G295));
  OAI21_X1  g447(.A(new_n871), .B1(G868), .B2(new_n820), .ZN(G331));
  XNOR2_X1  g448(.A(new_n824), .B(G286), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G301), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n874), .B(G171), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n862), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n878), .A3(new_n860), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT111), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n860), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(G37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT43), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(KEYINPUT44), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(G397));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n892));
  INV_X1    g467(.A(new_n500), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n492), .A2(new_n836), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n840), .A2(KEYINPUT108), .A3(new_n483), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n892), .B1(new_n896), .B2(G1384), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT112), .B(G40), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n472), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G1996), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n737), .B(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n793), .B(G2067), .Z(new_n904));
  OR2_X1    g479(.A1(new_n705), .A2(new_n707), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n705), .A2(new_n707), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(G1986), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n901), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT50), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT114), .B1(new_n896), .B2(G1384), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT114), .ZN(new_n912));
  INV_X1    g487(.A(G1384), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n842), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n910), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G1384), .B1(new_n492), .B2(new_n500), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n900), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n803), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT57), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n559), .A2(new_n920), .A3(new_n563), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n559), .B2(new_n563), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n892), .A2(G1384), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n894), .A2(new_n895), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n500), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n899), .B1(new_n916), .B2(KEYINPUT45), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT56), .B(G2072), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n919), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n911), .A2(new_n914), .A3(new_n910), .ZN(new_n933));
  INV_X1    g508(.A(new_n916), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n900), .B1(new_n934), .B2(KEYINPUT50), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1348), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n911), .A2(new_n914), .A3(new_n899), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n939), .A2(G2067), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n592), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n923), .B1(new_n919), .B2(new_n931), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n932), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n896), .A2(KEYINPUT114), .A3(G1384), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n912), .B1(new_n842), .B2(new_n913), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT50), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G1956), .B1(new_n946), .B2(new_n917), .ZN(new_n947));
  INV_X1    g522(.A(new_n931), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n947), .A2(new_n948), .B1(new_n922), .B2(new_n921), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT123), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n932), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT61), .B1(new_n942), .B2(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n938), .A2(new_n940), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT60), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n592), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n938), .A2(new_n940), .A3(KEYINPUT60), .A4(new_n593), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT58), .B(G1341), .Z(new_n961));
  NAND2_X1  g536(.A1(new_n939), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT121), .B(G1996), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n929), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n962), .A2(KEYINPUT122), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT122), .B1(new_n962), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n547), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT59), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT59), .B(new_n547), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n932), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n943), .B1(new_n960), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G1961), .B1(new_n933), .B2(new_n935), .ZN(new_n974));
  INV_X1    g549(.A(G2078), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT53), .B1(new_n929), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n978));
  XNOR2_X1  g553(.A(G171), .B(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G40), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(KEYINPUT53), .ZN(new_n981));
  NOR4_X1   g556(.A1(new_n927), .A2(new_n980), .A3(new_n472), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n982), .B2(new_n897), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n911), .B2(new_n914), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n899), .B1(G164), .B2(new_n925), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n985), .A2(new_n986), .A3(new_n981), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n987), .A2(new_n974), .A3(new_n976), .ZN(new_n988));
  INV_X1    g563(.A(new_n979), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(G303), .A2(G8), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT55), .Z(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n933), .A2(new_n993), .A3(new_n935), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n679), .B1(new_n927), .B2(new_n928), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n679), .C1(new_n927), .C2(new_n928), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(G8), .B(new_n992), .C1(new_n994), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n946), .A2(new_n993), .A3(new_n917), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n995), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n992), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n682), .A2(G1976), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n939), .A2(G8), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n939), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n570), .A2(new_n1012), .A3(new_n576), .ZN(new_n1013));
  INV_X1    g588(.A(G86), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n574), .B1(new_n523), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1015), .A2(KEYINPUT116), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(KEYINPUT116), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n573), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n1018), .B2(new_n1012), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1011), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n939), .A2(G8), .A3(new_n1005), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT119), .B1(new_n1010), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1008), .B(KEYINPUT115), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1011), .A2(new_n1020), .B1(new_n1022), .B2(KEYINPUT52), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n990), .B(new_n1004), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n911), .A2(new_n914), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n986), .B1(new_n1032), .B2(new_n892), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1033), .B2(G1966), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n933), .A2(new_n723), .A3(new_n935), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT120), .B(new_n757), .C1(new_n985), .C2(new_n986), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G286), .A2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1038), .B2(KEYINPUT124), .ZN(new_n1042));
  OAI211_X1 g617(.A(G8), .B(new_n1042), .C1(new_n1037), .C2(G286), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI211_X1 g619(.A(new_n1039), .B(new_n1042), .C1(new_n1037), .C2(G8), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n973), .A2(new_n1030), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1032), .A2(new_n892), .ZN(new_n1048));
  INV_X1    g623(.A(new_n986), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT120), .B1(new_n1050), .B2(new_n757), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1036), .A2(new_n1035), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(G168), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1010), .A2(new_n1024), .ZN(new_n1055));
  OAI21_X1  g630(.A(G8), .B1(new_n994), .B2(new_n999), .ZN(new_n1056));
  INV_X1    g631(.A(new_n992), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1000), .A2(KEYINPUT63), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1053), .B(new_n1004), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(KEYINPUT63), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n1011), .B(KEYINPUT117), .Z(new_n1063));
  XNOR2_X1  g638(.A(new_n1013), .B(KEYINPUT118), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G288), .A2(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1021), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1010), .A2(new_n1000), .A3(new_n1024), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1047), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1037), .A2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1042), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1038), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1043), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1071), .B1(new_n1075), .B2(new_n1040), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1040), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT62), .B(new_n1077), .C1(new_n1074), .C2(new_n1043), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1004), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n988), .A2(G301), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1076), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n909), .B1(new_n1070), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G290), .A2(G1986), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n901), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(KEYINPUT48), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(KEYINPUT48), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1087), .B(new_n1088), .C1(new_n901), .C2(new_n907), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT46), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n901), .A2(new_n902), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n904), .A2(new_n738), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1091), .B1(new_n1092), .B2(new_n901), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1091), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(KEYINPUT46), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1091), .A2(KEYINPUT125), .A3(new_n1090), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(new_n1098), .B(KEYINPUT47), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n903), .A2(new_n904), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1100), .A2(new_n906), .B1(G2067), .B2(new_n793), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1089), .B(new_n1099), .C1(new_n901), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1083), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT126), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1083), .A2(new_n1105), .A3(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g682(.A(G319), .ZN(new_n1109));
  NOR4_X1   g683(.A1(G229), .A2(G401), .A3(new_n1109), .A4(G227), .ZN(new_n1110));
  NAND3_X1  g684(.A1(new_n887), .A2(new_n856), .A3(new_n1110), .ZN(G225));
  INV_X1    g685(.A(G225), .ZN(G308));
endmodule


