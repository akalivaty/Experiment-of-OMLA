

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(n705), .ZN(n812) );
  XNOR2_X1 U555 ( .A(n751), .B(n520), .ZN(n519) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n520) );
  NOR2_X1 U557 ( .A1(n745), .A2(n744), .ZN(n750) );
  XNOR2_X1 U558 ( .A(n742), .B(KEYINPUT27), .ZN(n745) );
  INV_X1 U559 ( .A(G1384), .ZN(n521) );
  NAND2_X1 U560 ( .A1(n773), .A2(G286), .ZN(n767) );
  NAND2_X1 U561 ( .A1(n759), .A2(n760), .ZN(n773) );
  NAND2_X1 U562 ( .A1(n753), .A2(n519), .ZN(n755) );
  NAND2_X4 U563 ( .A1(n522), .A2(n521), .ZN(n705) );
  INV_X1 U564 ( .A(n704), .ZN(n522) );
  XNOR2_X2 U565 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n532) );
  BUF_X2 U566 ( .A(n921), .Z(n523) );
  NOR2_X1 U567 ( .A1(n535), .A2(n536), .ZN(n921) );
  NOR2_X2 U568 ( .A1(n775), .A2(n710), .ZN(n712) );
  AND2_X2 U569 ( .A1(n579), .A2(n578), .ZN(G160) );
  INV_X1 U570 ( .A(G2104), .ZN(n535) );
  INV_X1 U571 ( .A(KEYINPUT1), .ZN(n524) );
  OR2_X1 U572 ( .A1(n714), .A2(n706), .ZN(n707) );
  INV_X1 U573 ( .A(n616), .ZN(n741) );
  NAND2_X1 U574 ( .A1(G160), .A2(G40), .ZN(n811) );
  NOR2_X1 U575 ( .A1(n540), .A2(n539), .ZN(n704) );
  XNOR2_X1 U576 ( .A(n524), .B(n525), .ZN(n594) );
  BUF_X2 U577 ( .A(n574), .Z(n902) );
  NOR2_X2 U578 ( .A1(G543), .A2(G651), .ZN(n665) );
  XNOR2_X1 U579 ( .A(n605), .B(KEYINPUT15), .ZN(n616) );
  NAND2_X1 U580 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U581 ( .A(KEYINPUT70), .B(n548), .ZN(n525) );
  NOR2_X4 U582 ( .A1(n592), .A2(n591), .ZN(n1037) );
  BUF_X2 U583 ( .A(n594), .Z(n655) );
  INV_X1 U584 ( .A(KEYINPUT31), .ZN(n719) );
  INV_X1 U585 ( .A(n1052), .ZN(n797) );
  INV_X1 U586 ( .A(KEYINPUT30), .ZN(n711) );
  NOR2_X2 U587 ( .A1(n811), .A2(n705), .ZN(n714) );
  INV_X1 U588 ( .A(KEYINPUT64), .ZN(n787) );
  INV_X1 U589 ( .A(KEYINPUT102), .ZN(n780) );
  NOR2_X1 U590 ( .A1(n601), .A2(n600), .ZN(n604) );
  NOR2_X1 U591 ( .A1(n807), .A2(n530), .ZN(n808) );
  NOR2_X1 U592 ( .A1(G543), .A2(n547), .ZN(n548) );
  NOR2_X1 U593 ( .A1(n569), .A2(n568), .ZN(G171) );
  BUF_X1 U594 ( .A(n704), .Z(G164) );
  AND2_X1 U595 ( .A1(n1044), .A2(n857), .ZN(n526) );
  OR2_X1 U596 ( .A1(n741), .A2(n740), .ZN(n527) );
  NOR2_X1 U597 ( .A1(n802), .A2(n785), .ZN(n528) );
  AND2_X1 U598 ( .A1(KEYINPUT99), .A2(n1038), .ZN(n529) );
  AND2_X1 U599 ( .A1(n806), .A2(n805), .ZN(n530) );
  NOR2_X1 U600 ( .A1(n733), .A2(n529), .ZN(n734) );
  BUF_X1 U601 ( .A(n714), .Z(n743) );
  INV_X1 U602 ( .A(KEYINPUT29), .ZN(n754) );
  XNOR2_X1 U603 ( .A(n755), .B(n754), .ZN(n758) );
  INV_X1 U604 ( .A(KEYINPUT97), .ZN(n708) );
  INV_X1 U605 ( .A(KEYINPUT101), .ZN(n768) );
  INV_X1 U606 ( .A(n1045), .ZN(n785) );
  INV_X1 U607 ( .A(KEYINPUT105), .ZN(n795) );
  INV_X1 U608 ( .A(KEYINPUT80), .ZN(n598) );
  XNOR2_X1 U609 ( .A(n599), .B(n598), .ZN(n600) );
  NOR2_X1 U610 ( .A1(n659), .A2(G651), .ZN(n597) );
  NOR2_X1 U611 ( .A1(n842), .A2(n526), .ZN(n843) );
  BUF_X1 U612 ( .A(n616), .Z(n1034) );
  NAND2_X1 U613 ( .A1(n562), .A2(n561), .ZN(G299) );
  NOR2_X2 U614 ( .A1(n535), .A2(G2105), .ZN(n574) );
  NAND2_X1 U615 ( .A1(G102), .A2(n902), .ZN(n534) );
  NOR2_X1 U616 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XNOR2_X1 U617 ( .A(n532), .B(n531), .ZN(n624) );
  NAND2_X1 U618 ( .A1(G138), .A2(n624), .ZN(n533) );
  NAND2_X1 U619 ( .A1(n534), .A2(n533), .ZN(n540) );
  INV_X1 U620 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U621 ( .A1(G114), .A2(n523), .ZN(n538) );
  NOR2_X1 U622 ( .A1(G2104), .A2(n536), .ZN(n622) );
  NAND2_X1 U623 ( .A1(G126), .A2(n622), .ZN(n537) );
  NAND2_X1 U624 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U625 ( .A1(n665), .A2(G89), .ZN(n541) );
  XNOR2_X1 U626 ( .A(n541), .B(KEYINPUT4), .ZN(n544) );
  INV_X1 U627 ( .A(G651), .ZN(n547) );
  XOR2_X1 U628 ( .A(KEYINPUT0), .B(G543), .Z(n659) );
  OR2_X1 U629 ( .A1(n547), .A2(n659), .ZN(n542) );
  XNOR2_X1 U630 ( .A(KEYINPUT69), .B(n542), .ZN(n602) );
  BUF_X1 U631 ( .A(n602), .Z(n669) );
  NAND2_X1 U632 ( .A1(G76), .A2(n669), .ZN(n543) );
  NAND2_X1 U633 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U634 ( .A(KEYINPUT5), .B(n545), .ZN(n553) );
  BUF_X1 U635 ( .A(n597), .Z(n670) );
  NAND2_X1 U636 ( .A1(n670), .A2(G51), .ZN(n546) );
  XOR2_X1 U637 ( .A(KEYINPUT81), .B(n546), .Z(n550) );
  NAND2_X1 U638 ( .A1(G63), .A2(n655), .ZN(n549) );
  NAND2_X1 U639 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U640 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U641 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U642 ( .A(KEYINPUT7), .B(n554), .ZN(G168) );
  NAND2_X1 U643 ( .A1(G91), .A2(n665), .ZN(n555) );
  XNOR2_X1 U644 ( .A(n555), .B(KEYINPUT72), .ZN(n562) );
  NAND2_X1 U645 ( .A1(G53), .A2(n670), .ZN(n557) );
  NAND2_X1 U646 ( .A1(G78), .A2(n669), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U648 ( .A1(G65), .A2(n655), .ZN(n558) );
  XNOR2_X1 U649 ( .A(KEYINPUT73), .B(n558), .ZN(n559) );
  NOR2_X1 U650 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(n670), .A2(G52), .ZN(n564) );
  NAND2_X1 U653 ( .A1(G64), .A2(n655), .ZN(n563) );
  NAND2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U655 ( .A1(G90), .A2(n665), .ZN(n566) );
  NAND2_X1 U656 ( .A1(G77), .A2(n669), .ZN(n565) );
  NAND2_X1 U657 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U658 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  AND2_X1 U659 ( .A1(G452), .A2(G94), .ZN(G173) );
  AND2_X1 U660 ( .A1(G137), .A2(n624), .ZN(n573) );
  NAND2_X1 U661 ( .A1(G113), .A2(n523), .ZN(n571) );
  NAND2_X1 U662 ( .A1(G125), .A2(n622), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U664 ( .A1(n573), .A2(n572), .ZN(n579) );
  NAND2_X1 U665 ( .A1(G101), .A2(n574), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n575), .B(KEYINPUT23), .ZN(n577) );
  INV_X1 U667 ( .A(KEYINPUT66), .ZN(n576) );
  XNOR2_X1 U668 ( .A(n577), .B(n576), .ZN(n578) );
  INV_X1 U669 ( .A(G108), .ZN(G238) );
  INV_X1 U670 ( .A(G120), .ZN(G236) );
  INV_X1 U671 ( .A(G57), .ZN(G237) );
  INV_X1 U672 ( .A(G132), .ZN(G219) );
  NAND2_X1 U673 ( .A1(G7), .A2(G661), .ZN(n580) );
  XOR2_X1 U674 ( .A(n580), .B(KEYINPUT10), .Z(n862) );
  INV_X1 U675 ( .A(n862), .ZN(G223) );
  INV_X1 U676 ( .A(G567), .ZN(n698) );
  NOR2_X1 U677 ( .A1(n698), .A2(G223), .ZN(n581) );
  XNOR2_X1 U678 ( .A(n581), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U679 ( .A(G860), .B(KEYINPUT77), .Z(n611) );
  NAND2_X1 U680 ( .A1(G56), .A2(n655), .ZN(n582) );
  XNOR2_X1 U681 ( .A(n582), .B(KEYINPUT14), .ZN(n584) );
  NAND2_X1 U682 ( .A1(G43), .A2(n670), .ZN(n583) );
  NAND2_X1 U683 ( .A1(n584), .A2(n583), .ZN(n592) );
  XOR2_X1 U684 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n586) );
  NAND2_X1 U685 ( .A1(G81), .A2(n665), .ZN(n585) );
  XNOR2_X1 U686 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U687 ( .A(n587), .B(KEYINPUT75), .ZN(n589) );
  NAND2_X1 U688 ( .A1(n602), .A2(G68), .ZN(n588) );
  NAND2_X1 U689 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U690 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NAND2_X1 U691 ( .A1(n611), .A2(n1037), .ZN(n593) );
  XNOR2_X1 U692 ( .A(n593), .B(KEYINPUT78), .ZN(G153) );
  XNOR2_X1 U693 ( .A(G171), .B(KEYINPUT79), .ZN(G301) );
  NAND2_X1 U694 ( .A1(G868), .A2(G301), .ZN(n607) );
  NAND2_X1 U695 ( .A1(G92), .A2(n665), .ZN(n596) );
  NAND2_X1 U696 ( .A1(G66), .A2(n594), .ZN(n595) );
  NAND2_X1 U697 ( .A1(n596), .A2(n595), .ZN(n601) );
  NAND2_X1 U698 ( .A1(n597), .A2(G54), .ZN(n599) );
  NAND2_X1 U699 ( .A1(n602), .A2(G79), .ZN(n603) );
  INV_X1 U700 ( .A(G868), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n741), .A2(n614), .ZN(n606) );
  NAND2_X1 U702 ( .A1(n607), .A2(n606), .ZN(G284) );
  NOR2_X1 U703 ( .A1(G286), .A2(n614), .ZN(n609) );
  NOR2_X1 U704 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U705 ( .A1(n609), .A2(n608), .ZN(G297) );
  INV_X1 U706 ( .A(G559), .ZN(n610) );
  NOR2_X1 U707 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U708 ( .A1(n741), .A2(n612), .ZN(n613) );
  XOR2_X1 U709 ( .A(KEYINPUT16), .B(n613), .Z(G148) );
  NAND2_X1 U710 ( .A1(n1037), .A2(n614), .ZN(n615) );
  XOR2_X1 U711 ( .A(KEYINPUT82), .B(n615), .Z(n619) );
  NAND2_X1 U712 ( .A1(G868), .A2(n1034), .ZN(n617) );
  NOR2_X1 U713 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U714 ( .A1(n619), .A2(n618), .ZN(G282) );
  XOR2_X1 U715 ( .A(G2100), .B(KEYINPUT84), .Z(n632) );
  NAND2_X1 U716 ( .A1(G99), .A2(n902), .ZN(n621) );
  NAND2_X1 U717 ( .A1(G111), .A2(n523), .ZN(n620) );
  NAND2_X1 U718 ( .A1(n621), .A2(n620), .ZN(n630) );
  BUF_X1 U719 ( .A(n622), .Z(n922) );
  NAND2_X1 U720 ( .A1(n922), .A2(G123), .ZN(n623) );
  XNOR2_X1 U721 ( .A(n623), .B(KEYINPUT18), .ZN(n627) );
  BUF_X1 U722 ( .A(n624), .Z(n625) );
  NAND2_X1 U723 ( .A1(G135), .A2(n625), .ZN(n626) );
  NAND2_X1 U724 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U725 ( .A(KEYINPUT83), .B(n628), .Z(n629) );
  NOR2_X1 U726 ( .A1(n630), .A2(n629), .ZN(n1023) );
  XNOR2_X1 U727 ( .A(n1023), .B(G2096), .ZN(n631) );
  NAND2_X1 U728 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U729 ( .A1(n670), .A2(G55), .ZN(n634) );
  NAND2_X1 U730 ( .A1(G67), .A2(n655), .ZN(n633) );
  NAND2_X1 U731 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U732 ( .A1(G93), .A2(n665), .ZN(n636) );
  NAND2_X1 U733 ( .A1(G80), .A2(n669), .ZN(n635) );
  NAND2_X1 U734 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U735 ( .A1(n638), .A2(n637), .ZN(n684) );
  NAND2_X1 U736 ( .A1(G559), .A2(n1034), .ZN(n639) );
  XOR2_X1 U737 ( .A(n639), .B(n1037), .Z(n682) );
  NOR2_X1 U738 ( .A1(G860), .A2(n682), .ZN(n640) );
  XOR2_X1 U739 ( .A(KEYINPUT85), .B(n640), .Z(n641) );
  XNOR2_X1 U740 ( .A(n684), .B(n641), .ZN(G145) );
  NAND2_X1 U741 ( .A1(n655), .A2(G62), .ZN(n642) );
  XNOR2_X1 U742 ( .A(n642), .B(KEYINPUT87), .ZN(n649) );
  NAND2_X1 U743 ( .A1(G88), .A2(n665), .ZN(n644) );
  NAND2_X1 U744 ( .A1(G75), .A2(n669), .ZN(n643) );
  NAND2_X1 U745 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U746 ( .A(KEYINPUT88), .B(n645), .Z(n647) );
  NAND2_X1 U747 ( .A1(n670), .A2(G50), .ZN(n646) );
  NAND2_X1 U748 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U749 ( .A1(n649), .A2(n648), .ZN(G166) );
  INV_X1 U750 ( .A(G166), .ZN(G303) );
  NAND2_X1 U751 ( .A1(G86), .A2(n665), .ZN(n651) );
  NAND2_X1 U752 ( .A1(G48), .A2(n670), .ZN(n650) );
  NAND2_X1 U753 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U754 ( .A1(n669), .A2(G73), .ZN(n652) );
  XOR2_X1 U755 ( .A(KEYINPUT2), .B(n652), .Z(n653) );
  NOR2_X1 U756 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U757 ( .A1(G61), .A2(n655), .ZN(n656) );
  NAND2_X1 U758 ( .A1(n657), .A2(n656), .ZN(G305) );
  NAND2_X1 U759 ( .A1(G74), .A2(G651), .ZN(n658) );
  XNOR2_X1 U760 ( .A(n658), .B(KEYINPUT86), .ZN(n664) );
  NAND2_X1 U761 ( .A1(G49), .A2(n670), .ZN(n661) );
  NAND2_X1 U762 ( .A1(G87), .A2(n659), .ZN(n660) );
  NAND2_X1 U763 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U764 ( .A1(n594), .A2(n662), .ZN(n663) );
  NAND2_X1 U765 ( .A1(n664), .A2(n663), .ZN(G288) );
  NAND2_X1 U766 ( .A1(n665), .A2(G85), .ZN(n666) );
  XNOR2_X1 U767 ( .A(KEYINPUT68), .B(n666), .ZN(n668) );
  NAND2_X1 U768 ( .A1(G60), .A2(n594), .ZN(n667) );
  NAND2_X1 U769 ( .A1(n668), .A2(n667), .ZN(n674) );
  NAND2_X1 U770 ( .A1(n669), .A2(G72), .ZN(n672) );
  NAND2_X1 U771 ( .A1(n670), .A2(G47), .ZN(n671) );
  NAND2_X1 U772 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U773 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U774 ( .A(KEYINPUT71), .B(n675), .ZN(G290) );
  XOR2_X1 U775 ( .A(G299), .B(n684), .Z(n680) );
  XOR2_X1 U776 ( .A(G303), .B(G305), .Z(n678) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(KEYINPUT19), .ZN(n676) );
  XNOR2_X1 U778 ( .A(n676), .B(G288), .ZN(n677) );
  XNOR2_X1 U779 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U780 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U781 ( .A(n681), .B(G290), .ZN(n935) );
  XOR2_X1 U782 ( .A(n682), .B(n935), .Z(n683) );
  NAND2_X1 U783 ( .A1(n683), .A2(G868), .ZN(n686) );
  OR2_X1 U784 ( .A1(G868), .A2(n684), .ZN(n685) );
  NAND2_X1 U785 ( .A1(n686), .A2(n685), .ZN(G295) );
  NAND2_X1 U786 ( .A1(G2084), .A2(G2078), .ZN(n688) );
  XOR2_X1 U787 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n687) );
  XNOR2_X1 U788 ( .A(n688), .B(n687), .ZN(n689) );
  NAND2_X1 U789 ( .A1(G2090), .A2(n689), .ZN(n690) );
  XNOR2_X1 U790 ( .A(KEYINPUT21), .B(n690), .ZN(n691) );
  NAND2_X1 U791 ( .A1(n691), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U792 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U793 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  NOR2_X1 U794 ( .A1(G220), .A2(G219), .ZN(n692) );
  XOR2_X1 U795 ( .A(KEYINPUT22), .B(n692), .Z(n693) );
  NOR2_X1 U796 ( .A1(G218), .A2(n693), .ZN(n694) );
  NAND2_X1 U797 ( .A1(G96), .A2(n694), .ZN(n868) );
  NAND2_X1 U798 ( .A1(G2106), .A2(n868), .ZN(n695) );
  XNOR2_X1 U799 ( .A(n695), .B(KEYINPUT91), .ZN(n700) );
  NOR2_X1 U800 ( .A1(G236), .A2(G238), .ZN(n696) );
  NAND2_X1 U801 ( .A1(G69), .A2(n696), .ZN(n697) );
  NOR2_X1 U802 ( .A1(G237), .A2(n697), .ZN(n867) );
  NOR2_X1 U803 ( .A1(n698), .A2(n867), .ZN(n699) );
  NOR2_X1 U804 ( .A1(n700), .A2(n699), .ZN(G319) );
  INV_X1 U805 ( .A(G319), .ZN(n702) );
  NAND2_X1 U806 ( .A1(G483), .A2(G661), .ZN(n701) );
  NOR2_X1 U807 ( .A1(n702), .A2(n701), .ZN(n866) );
  NAND2_X1 U808 ( .A1(n866), .A2(G36), .ZN(G176) );
  INV_X1 U809 ( .A(G8), .ZN(n706) );
  XNOR2_X1 U810 ( .A(n707), .B(KEYINPUT96), .ZN(n761) );
  NOR2_X1 U811 ( .A1(n761), .A2(G1966), .ZN(n709) );
  XNOR2_X1 U812 ( .A(n709), .B(n708), .ZN(n775) );
  INV_X1 U813 ( .A(n714), .ZN(n762) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n762), .ZN(n772) );
  OR2_X1 U815 ( .A1(n706), .A2(n772), .ZN(n710) );
  XNOR2_X1 U816 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U817 ( .A1(n713), .A2(G168), .ZN(n718) );
  XOR2_X1 U818 ( .A(G1961), .B(KEYINPUT98), .Z(n956) );
  NAND2_X1 U819 ( .A1(n956), .A2(n762), .ZN(n716) );
  XNOR2_X1 U820 ( .A(G2078), .B(KEYINPUT25), .ZN(n991) );
  NAND2_X1 U821 ( .A1(n743), .A2(n991), .ZN(n715) );
  NAND2_X1 U822 ( .A1(n716), .A2(n715), .ZN(n756) );
  NOR2_X1 U823 ( .A1(G171), .A2(n756), .ZN(n717) );
  NOR2_X1 U824 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U825 ( .A(n720), .B(n719), .ZN(n760) );
  XOR2_X1 U826 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n726) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n726), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n741), .A2(G2067), .ZN(n722) );
  NAND2_X1 U829 ( .A1(G1996), .A2(n726), .ZN(n721) );
  NAND2_X1 U830 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U831 ( .A1(KEYINPUT99), .A2(n723), .ZN(n724) );
  NOR2_X1 U832 ( .A1(n762), .A2(n724), .ZN(n725) );
  INV_X1 U833 ( .A(n725), .ZN(n735) );
  NAND2_X1 U834 ( .A1(G1348), .A2(n741), .ZN(n730) );
  INV_X1 U835 ( .A(n726), .ZN(n728) );
  INV_X1 U836 ( .A(G1341), .ZN(n1038) );
  NOR2_X1 U837 ( .A1(KEYINPUT99), .A2(n1038), .ZN(n727) );
  NOR2_X1 U838 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U839 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U840 ( .A1(n731), .A2(n762), .ZN(n732) );
  NAND2_X1 U841 ( .A1(n732), .A2(n1037), .ZN(n733) );
  NAND2_X1 U842 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U843 ( .A1(n737), .A2(n736), .ZN(n748) );
  NAND2_X1 U844 ( .A1(G1348), .A2(n762), .ZN(n739) );
  NAND2_X1 U845 ( .A1(G2067), .A2(n743), .ZN(n738) );
  NAND2_X1 U846 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U847 ( .A1(n743), .A2(G2072), .ZN(n742) );
  INV_X1 U848 ( .A(G1956), .ZN(n870) );
  NOR2_X1 U849 ( .A1(n870), .A2(n743), .ZN(n744) );
  INV_X1 U850 ( .A(G299), .ZN(n749) );
  NAND2_X1 U851 ( .A1(n750), .A2(n749), .ZN(n746) );
  NAND2_X1 U852 ( .A1(n527), .A2(n746), .ZN(n747) );
  OR2_X1 U853 ( .A1(n748), .A2(n747), .ZN(n753) );
  NOR2_X1 U854 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U855 ( .A1(n756), .A2(G171), .ZN(n757) );
  NAND2_X1 U856 ( .A1(n758), .A2(n757), .ZN(n759) );
  BUF_X1 U857 ( .A(n761), .Z(n802) );
  NOR2_X1 U858 ( .A1(n802), .A2(G1971), .ZN(n764) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n765), .A2(G303), .ZN(n766) );
  NAND2_X1 U862 ( .A1(n767), .A2(n766), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n770), .A2(G8), .ZN(n771) );
  XNOR2_X1 U865 ( .A(n771), .B(KEYINPUT32), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G8), .A2(n772), .ZN(n777) );
  XOR2_X1 U867 ( .A(KEYINPUT100), .B(n773), .Z(n774) );
  NOR2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n781) );
  XNOR2_X1 U871 ( .A(n781), .B(n780), .ZN(n799) );
  INV_X1 U872 ( .A(n799), .ZN(n783) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n790) );
  NOR2_X1 U874 ( .A1(G1971), .A2(G303), .ZN(n782) );
  NOR2_X1 U875 ( .A1(n790), .A2(n782), .ZN(n1041) );
  NAND2_X1 U876 ( .A1(n783), .A2(n1041), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G288), .A2(G1976), .ZN(n784) );
  XOR2_X1 U878 ( .A(KEYINPUT103), .B(n784), .Z(n1045) );
  NAND2_X1 U879 ( .A1(n786), .A2(n528), .ZN(n788) );
  XNOR2_X1 U880 ( .A(n788), .B(n787), .ZN(n789) );
  NOR2_X1 U881 ( .A1(n789), .A2(KEYINPUT33), .ZN(n794) );
  NAND2_X1 U882 ( .A1(KEYINPUT33), .A2(n790), .ZN(n791) );
  NOR2_X1 U883 ( .A1(n802), .A2(n791), .ZN(n792) );
  XNOR2_X1 U884 ( .A(n792), .B(KEYINPUT104), .ZN(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n796) );
  XNOR2_X1 U886 ( .A(n796), .B(n795), .ZN(n798) );
  XNOR2_X1 U887 ( .A(G1981), .B(G305), .ZN(n1052) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n809) );
  NAND2_X1 U889 ( .A1(G166), .A2(G8), .ZN(n800) );
  NOR2_X1 U890 ( .A1(G2090), .A2(n800), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n799), .A2(n801), .ZN(n803) );
  INV_X1 U892 ( .A(n802), .ZN(n805) );
  NOR2_X1 U893 ( .A1(n803), .A2(n805), .ZN(n807) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n804), .B(KEYINPUT24), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(KEYINPUT106), .ZN(n844) );
  NOR2_X1 U898 ( .A1(n812), .A2(n811), .ZN(n857) );
  XNOR2_X1 U899 ( .A(G2067), .B(KEYINPUT37), .ZN(n845) );
  NAND2_X1 U900 ( .A1(G104), .A2(n902), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G140), .A2(n625), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U903 ( .A(KEYINPUT34), .B(n815), .ZN(n820) );
  NAND2_X1 U904 ( .A1(G116), .A2(n523), .ZN(n817) );
  NAND2_X1 U905 ( .A1(G128), .A2(n922), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  XOR2_X1 U907 ( .A(KEYINPUT35), .B(n818), .Z(n819) );
  NOR2_X1 U908 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U909 ( .A(KEYINPUT36), .B(n821), .ZN(n899) );
  NOR2_X1 U910 ( .A1(n845), .A2(n899), .ZN(n1020) );
  NAND2_X1 U911 ( .A1(n857), .A2(n1020), .ZN(n854) );
  NAND2_X1 U912 ( .A1(n523), .A2(G117), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(KEYINPUT92), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G129), .A2(n922), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G105), .A2(n902), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT93), .ZN(n826) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT38), .ZN(n827) );
  NOR2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U920 ( .A(n829), .B(KEYINPUT94), .ZN(n831) );
  NAND2_X1 U921 ( .A1(G141), .A2(n625), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n900) );
  NAND2_X1 U923 ( .A1(G1996), .A2(n900), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT95), .ZN(n840) );
  INV_X1 U925 ( .A(G1991), .ZN(n982) );
  NAND2_X1 U926 ( .A1(G95), .A2(n902), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G131), .A2(n625), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n838) );
  NAND2_X1 U929 ( .A1(G107), .A2(n523), .ZN(n836) );
  NAND2_X1 U930 ( .A1(G119), .A2(n922), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n918) );
  NOR2_X1 U933 ( .A1(n982), .A2(n918), .ZN(n839) );
  NOR2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n1018) );
  INV_X1 U935 ( .A(n1018), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n841), .A2(n857), .ZN(n846) );
  NAND2_X1 U937 ( .A1(n854), .A2(n846), .ZN(n842) );
  XNOR2_X1 U938 ( .A(G1986), .B(G290), .ZN(n1044) );
  NAND2_X1 U939 ( .A1(n844), .A2(n843), .ZN(n860) );
  NAND2_X1 U940 ( .A1(n845), .A2(n899), .ZN(n1010) );
  NOR2_X1 U941 ( .A1(G1996), .A2(n900), .ZN(n1013) );
  INV_X1 U942 ( .A(n846), .ZN(n850) );
  AND2_X1 U943 ( .A1(n982), .A2(n918), .ZN(n1019) );
  NOR2_X1 U944 ( .A1(G1986), .A2(G290), .ZN(n847) );
  XOR2_X1 U945 ( .A(n847), .B(KEYINPUT107), .Z(n848) );
  NOR2_X1 U946 ( .A1(n1019), .A2(n848), .ZN(n849) );
  NOR2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U948 ( .A1(n1013), .A2(n851), .ZN(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT39), .B(n852), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n853), .B(KEYINPUT108), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n1010), .A2(n856), .ZN(n858) );
  NAND2_X1 U953 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U954 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U955 ( .A(n861), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U956 ( .A1(G2106), .A2(n862), .ZN(G217) );
  AND2_X1 U957 ( .A1(G15), .A2(G2), .ZN(n863) );
  NAND2_X1 U958 ( .A1(G661), .A2(n863), .ZN(G259) );
  NAND2_X1 U959 ( .A1(G3), .A2(G1), .ZN(n864) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(n864), .Z(n865) );
  NAND2_X1 U961 ( .A1(n866), .A2(n865), .ZN(G188) );
  INV_X1 U963 ( .A(G96), .ZN(G221) );
  INV_X1 U964 ( .A(n867), .ZN(n869) );
  NOR2_X1 U965 ( .A1(n869), .A2(n868), .ZN(G325) );
  INV_X1 U966 ( .A(G325), .ZN(G261) );
  XOR2_X1 U967 ( .A(KEYINPUT41), .B(G1976), .Z(n872) );
  XOR2_X1 U968 ( .A(G1961), .B(n870), .Z(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U970 ( .A(n873), .B(KEYINPUT112), .Z(n875) );
  XOR2_X1 U971 ( .A(G1996), .B(n982), .Z(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U973 ( .A(G1971), .B(G1966), .Z(n877) );
  XNOR2_X1 U974 ( .A(G1986), .B(G1981), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U976 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U977 ( .A(KEYINPUT111), .B(G2474), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(G229) );
  XOR2_X1 U979 ( .A(G2100), .B(KEYINPUT43), .Z(n883) );
  XNOR2_X1 U980 ( .A(G2090), .B(G2678), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(n884), .B(KEYINPUT110), .Z(n886) );
  XNOR2_X1 U983 ( .A(G2067), .B(G2072), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U985 ( .A(KEYINPUT42), .B(G2096), .Z(n888) );
  XNOR2_X1 U986 ( .A(G2084), .B(G2078), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(G227) );
  NAND2_X1 U989 ( .A1(G124), .A2(n922), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n891), .B(KEYINPUT44), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G136), .A2(n625), .ZN(n892) );
  XOR2_X1 U992 ( .A(KEYINPUT113), .B(n892), .Z(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n898) );
  NAND2_X1 U994 ( .A1(G100), .A2(n902), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G112), .A2(n523), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(G162) );
  XNOR2_X1 U998 ( .A(n1023), .B(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n914) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n902), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n625), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n523), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(G127), .A2(n922), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1006 ( .A(KEYINPUT116), .B(n907), .Z(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT47), .B(n908), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n1006) );
  XOR2_X1 U1009 ( .A(n1006), .B(G162), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G164), .B(G160), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1012 ( .A(n914), .B(n913), .Z(n920) );
  XOR2_X1 U1013 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n916) );
  XNOR2_X1 U1014 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n933) );
  NAND2_X1 U1018 ( .A1(G118), .A2(n523), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(G130), .A2(n922), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n931) );
  NAND2_X1 U1021 ( .A1(n902), .A2(G106), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT114), .B(n925), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n625), .A2(G142), .ZN(n926) );
  XOR2_X1 U1024 ( .A(KEYINPUT115), .B(n926), .Z(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1026 ( .A(n929), .B(KEYINPUT45), .Z(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(n933), .B(n932), .Z(n934) );
  NOR2_X1 U1029 ( .A1(G37), .A2(n934), .ZN(G395) );
  XOR2_X1 U1030 ( .A(KEYINPUT119), .B(n1034), .Z(n936) );
  XOR2_X1 U1031 ( .A(n936), .B(n935), .Z(n938) );
  XNOR2_X1 U1032 ( .A(G171), .B(n1037), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n938), .B(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(G286), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(G37), .A2(n940), .ZN(G397) );
  XOR2_X1 U1036 ( .A(G2451), .B(G2430), .Z(n942) );
  XNOR2_X1 U1037 ( .A(G2438), .B(G2443), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(n942), .B(n941), .ZN(n948) );
  XOR2_X1 U1039 ( .A(G2435), .B(G2454), .Z(n944) );
  XOR2_X1 U1040 ( .A(G1348), .B(n1038), .Z(n943) );
  XNOR2_X1 U1041 ( .A(n944), .B(n943), .ZN(n946) );
  XOR2_X1 U1042 ( .A(G2446), .B(G2427), .Z(n945) );
  XNOR2_X1 U1043 ( .A(n946), .B(n945), .ZN(n947) );
  XOR2_X1 U1044 ( .A(n948), .B(n947), .Z(n949) );
  NAND2_X1 U1045 ( .A1(G14), .A2(n949), .ZN(n955) );
  NAND2_X1 U1046 ( .A1(G319), .A2(n955), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(G229), .A2(G227), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(KEYINPUT49), .B(n950), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(G395), .A2(G397), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(G225) );
  INV_X1 U1052 ( .A(G225), .ZN(G308) );
  INV_X1 U1053 ( .A(G69), .ZN(G235) );
  INV_X1 U1054 ( .A(n955), .ZN(G401) );
  XNOR2_X1 U1055 ( .A(n956), .B(G5), .ZN(n978) );
  XOR2_X1 U1056 ( .A(G1966), .B(G21), .Z(n965) );
  XOR2_X1 U1057 ( .A(G1976), .B(G23), .Z(n959) );
  XOR2_X1 U1058 ( .A(KEYINPUT126), .B(G24), .Z(n957) );
  XNOR2_X1 U1059 ( .A(n957), .B(G1986), .ZN(n958) );
  NAND2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1061 ( .A(KEYINPUT125), .B(G1971), .Z(n960) );
  XNOR2_X1 U1062 ( .A(G22), .B(n960), .ZN(n961) );
  NOR2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n976) );
  XOR2_X1 U1066 ( .A(G20), .B(G1956), .Z(n969) );
  XNOR2_X1 U1067 ( .A(G1981), .B(G6), .ZN(n967) );
  XOR2_X1 U1068 ( .A(G19), .B(n1038), .Z(n966) );
  NOR2_X1 U1069 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1071 ( .A(KEYINPUT59), .B(G1348), .Z(n970) );
  XNOR2_X1 U1072 ( .A(G4), .B(n970), .ZN(n971) );
  NOR2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1074 ( .A(KEYINPUT60), .B(n973), .Z(n974) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(n974), .ZN(n975) );
  NOR2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1078 ( .A(n979), .B(KEYINPUT127), .ZN(n980) );
  XOR2_X1 U1079 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1080 ( .A1(G16), .A2(n981), .ZN(n1005) );
  XNOR2_X1 U1081 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n1029) );
  XNOR2_X1 U1082 ( .A(G2090), .B(G35), .ZN(n996) );
  XOR2_X1 U1083 ( .A(n982), .B(G25), .Z(n984) );
  XNOR2_X1 U1084 ( .A(G33), .B(G2072), .ZN(n983) );
  NOR2_X1 U1085 ( .A1(n984), .A2(n983), .ZN(n990) );
  XOR2_X1 U1086 ( .A(G1996), .B(G32), .Z(n985) );
  NAND2_X1 U1087 ( .A1(n985), .A2(G28), .ZN(n988) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(G2067), .ZN(n986) );
  XNOR2_X1 U1089 ( .A(G26), .B(n986), .ZN(n987) );
  NOR2_X1 U1090 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1091 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1092 ( .A(G27), .B(n991), .Z(n992) );
  NOR2_X1 U1093 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1094 ( .A(KEYINPUT53), .B(n994), .ZN(n995) );
  NOR2_X1 U1095 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1096 ( .A(G2084), .B(G34), .Z(n997) );
  XNOR2_X1 U1097 ( .A(KEYINPUT54), .B(n997), .ZN(n998) );
  NAND2_X1 U1098 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1099 ( .A(n1029), .B(n1000), .ZN(n1002) );
  INV_X1 U1100 ( .A(G29), .ZN(n1001) );
  NAND2_X1 U1101 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1003), .ZN(n1004) );
  NOR2_X1 U1103 ( .A1(n1005), .A2(n1004), .ZN(n1033) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1006), .Z(n1008) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1007) );
  NOR2_X1 U1106 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1107 ( .A(n1009), .B(KEYINPUT50), .ZN(n1011) );
  NAND2_X1 U1108 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1109 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1110 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1111 ( .A(n1014), .B(KEYINPUT51), .ZN(n1015) );
  NOR2_X1 U1112 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1113 ( .A1(n1018), .A2(n1017), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(G160), .B(G2084), .ZN(n1022) );
  NOR2_X1 U1115 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1116 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NOR2_X1 U1117 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1118 ( .A(KEYINPUT120), .B(n1025), .Z(n1026) );
  NOR2_X1 U1119 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1120 ( .A(KEYINPUT52), .B(n1028), .ZN(n1030) );
  NAND2_X1 U1121 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1122 ( .A1(n1031), .A2(G29), .ZN(n1032) );
  NAND2_X1 U1123 ( .A1(n1033), .A2(n1032), .ZN(n1060) );
  XOR2_X1 U1124 ( .A(G171), .B(G1961), .Z(n1036) );
  XOR2_X1 U1125 ( .A(n1034), .B(G1348), .Z(n1035) );
  NOR2_X1 U1126 ( .A1(n1036), .A2(n1035), .ZN(n1050) );
  XOR2_X1 U1127 ( .A(n1038), .B(n1037), .Z(n1040) );
  NAND2_X1 U1128 ( .A1(G1971), .A2(G303), .ZN(n1039) );
  NAND2_X1 U1129 ( .A1(n1040), .A2(n1039), .ZN(n1048) );
  XOR2_X1 U1130 ( .A(G299), .B(G1956), .Z(n1042) );
  NAND2_X1 U1131 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NOR2_X1 U1132 ( .A1(n1044), .A2(n1043), .ZN(n1046) );
  NAND2_X1 U1133 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1134 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NAND2_X1 U1135 ( .A1(n1050), .A2(n1049), .ZN(n1056) );
  XNOR2_X1 U1136 ( .A(G1966), .B(G168), .ZN(n1051) );
  XNOR2_X1 U1137 ( .A(n1051), .B(KEYINPUT123), .ZN(n1053) );
  NOR2_X1 U1138 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  XNOR2_X1 U1139 ( .A(KEYINPUT57), .B(n1054), .ZN(n1055) );
  NOR2_X1 U1140 ( .A1(n1056), .A2(n1055), .ZN(n1058) );
  XOR2_X1 U1141 ( .A(KEYINPUT56), .B(G16), .Z(n1057) );
  NOR2_X1 U1142 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  NOR2_X1 U1143 ( .A1(n1060), .A2(n1059), .ZN(n1061) );
  XOR2_X1 U1144 ( .A(n1061), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1145 ( .A(G150), .ZN(G311) );
endmodule

