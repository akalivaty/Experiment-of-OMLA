//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n465), .A2(G136), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT66), .Z(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n466), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n484), .B(new_n486), .C1(new_n463), .C2(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n466), .A2(G138), .ZN(new_n488));
  OR2_X1    g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n494), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n500), .B2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(KEYINPUT69), .B2(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(G88), .B1(G50), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n505), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n513), .A2(G51), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT71), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n504), .A2(new_n501), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n526), .A2(new_n527), .A3(new_n502), .A4(new_n523), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n522), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(KEYINPUT72), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n526), .A2(G89), .A3(new_n509), .A4(new_n502), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n531), .A2(KEYINPUT73), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  AOI211_X1 g114(.A(new_n539), .B(new_n522), .C1(new_n525), .C2(new_n528), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n530), .A2(new_n538), .A3(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n511), .A2(G90), .ZN(new_n542));
  INV_X1    g117(.A(new_n513), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT74), .B(G52), .Z(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n526), .A2(G64), .A3(new_n502), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  XNOR2_X1  g125(.A(KEYINPUT75), .B(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n511), .A2(G81), .B1(new_n513), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n505), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n513), .A2(G53), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n513), .A2(new_n566), .A3(G53), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n511), .A2(G91), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n526), .A2(G65), .A3(new_n502), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  OR2_X1    g148(.A1(new_n545), .A2(new_n549), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  NAND4_X1  g150(.A1(new_n526), .A2(G87), .A3(new_n509), .A4(new_n502), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n513), .A2(G49), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n546), .B1(new_n505), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(KEYINPUT76), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n577), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n580), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n511), .A2(G86), .B1(G48), .B2(new_n513), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n505), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n505), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n513), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n511), .A2(G85), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G290));
  NAND4_X1  g175(.A1(new_n526), .A2(G92), .A3(new_n509), .A4(new_n502), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n505), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n543), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n513), .A2(KEYINPUT77), .ZN(new_n610));
  AOI22_X1  g185(.A1(G651), .A2(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G171), .ZN(G284));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G171), .ZN(G321));
  NAND2_X1  g191(.A1(G299), .A2(new_n613), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n613), .ZN(G280));
  XOR2_X1   g193(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g194(.A(new_n612), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT79), .B(G559), .Z(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(G860), .B2(new_n621), .ZN(G148));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n623));
  INV_X1    g198(.A(new_n621), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n612), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n603), .A2(KEYINPUT80), .A3(new_n611), .A4(new_n621), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  MUX2_X1   g202(.A(new_n557), .B(new_n627), .S(G868), .Z(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(new_n464), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n467), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2100), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n465), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n477), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n466), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT81), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n634), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2430), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n648), .A2(KEYINPUT83), .A3(KEYINPUT14), .ZN(new_n649));
  AOI21_X1  g224(.A(KEYINPUT83), .B1(new_n648), .B2(KEYINPUT14), .ZN(new_n650));
  OAI22_X1  g225(.A1(new_n649), .A2(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT17), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n666), .B2(new_n664), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT84), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n666), .A3(new_n664), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n666), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n665), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n690), .B(new_n689), .S(new_n682), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT85), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT86), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(new_n698), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT87), .B(G1986), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n699), .B2(new_n700), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(G229));
  NOR2_X1   g281(.A1(G29), .A2(G35), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G162), .B2(G29), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G2090), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT94), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G21), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G168), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1966), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(G19), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n558), .B2(new_n712), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT91), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1341), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2078), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n712), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n712), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1961), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n722), .A2(G33), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n465), .A2(G139), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n630), .A2(G127), .ZN(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n466), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n730), .B1(new_n740), .B2(new_n722), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2072), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT30), .B(G28), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n743), .A2(new_n722), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n641), .B2(new_n722), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G4), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n620), .B2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G1348), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n722), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  OAI211_X1 g328(.A(G140), .B(new_n466), .C1(new_n462), .C2(new_n463), .ZN(new_n754));
  OAI211_X1 g329(.A(G128), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n755));
  INV_X1    g330(.A(G116), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G104), .C2(G2105), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n754), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n722), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n473), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2084), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n748), .A2(new_n751), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  NOR4_X1   g344(.A1(new_n721), .A2(new_n726), .A3(new_n729), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n709), .A2(G2090), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n712), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT95), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT96), .B(G1956), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n722), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n465), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n477), .A2(G129), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n467), .A2(G105), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT26), .Z(new_n783));
  NAND4_X1  g358(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n722), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G1348), .B2(new_n750), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n771), .A2(new_n777), .A3(new_n789), .ZN(new_n790));
  AND4_X1   g365(.A1(new_n711), .A2(new_n716), .A3(new_n770), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n712), .A2(G24), .ZN(new_n792));
  AND3_X1   g367(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n712), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1986), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n722), .A2(G25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n465), .A2(G131), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n477), .A2(G119), .ZN(new_n798));
  OR2_X1    g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n722), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n712), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n712), .ZN(new_n810));
  INV_X1    g385(.A(G1971), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n712), .A2(G23), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n584), .A2(new_n580), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n712), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT33), .B(G1976), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n808), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n795), .B(new_n805), .C1(new_n818), .C2(KEYINPUT34), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT88), .Z(new_n820));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n818), .B2(KEYINPUT34), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(KEYINPUT36), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n791), .A2(new_n823), .A3(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n557), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n505), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G651), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n513), .A2(G55), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n511), .A2(G93), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n556), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n830), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n557), .A2(new_n837), .A3(new_n829), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT38), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n620), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT98), .B(G860), .Z(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n838), .A2(new_n848), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  NAND2_X1  g427(.A1(new_n465), .A2(G142), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n477), .A2(G130), .ZN(new_n854));
  OR2_X1    g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n740), .ZN(new_n859));
  INV_X1    g434(.A(new_n785), .ZN(new_n860));
  INV_X1    g435(.A(new_n498), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n487), .B(KEYINPUT99), .C1(new_n491), .C2(new_n492), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n484), .B1(new_n462), .B2(new_n463), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT4), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT68), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n486), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT99), .B1(new_n868), .B2(new_n487), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n861), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n759), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n493), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n862), .ZN(new_n874));
  INV_X1    g449(.A(new_n759), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n861), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(KEYINPUT100), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT100), .B1(new_n871), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n875), .B1(new_n874), .B2(new_n861), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n498), .B(new_n759), .C1(new_n873), .C2(new_n862), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(KEYINPUT100), .A3(new_n876), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n785), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n859), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n784), .B1(new_n881), .B2(new_n882), .ZN(new_n887));
  INV_X1    g462(.A(new_n784), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n871), .A2(new_n888), .A3(new_n876), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n859), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n858), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n632), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n883), .A2(new_n785), .A3(new_n884), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n785), .B1(new_n883), .B2(new_n884), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n740), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n890), .A3(new_n857), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n892), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n893), .B1(new_n892), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n801), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n640), .B(G160), .ZN(new_n901));
  XNOR2_X1  g476(.A(G162), .B(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n886), .A2(new_n858), .A3(new_n891), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n857), .B1(new_n896), .B2(new_n890), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n632), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n892), .A2(new_n897), .A3(new_n893), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n802), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT101), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n900), .A2(new_n907), .A3(new_n910), .A4(new_n902), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n902), .B1(new_n900), .B2(new_n907), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(G37), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n625), .A2(KEYINPUT102), .A3(new_n626), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT102), .B1(new_n625), .B2(new_n626), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n842), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n627), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n842), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n625), .A2(KEYINPUT102), .A3(new_n626), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n565), .A2(new_n567), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n526), .A2(G91), .A3(new_n509), .A4(new_n502), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n546), .B1(new_n569), .B2(new_n570), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT103), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n568), .A2(new_n572), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n931), .A2(new_n933), .A3(new_n603), .A4(new_n611), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n612), .A2(KEYINPUT103), .A3(G299), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT41), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT41), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n921), .A2(new_n926), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n935), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n921), .B2(new_n926), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT105), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n919), .A2(new_n920), .A3(new_n842), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n924), .B1(new_n923), .B2(new_n925), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n921), .A2(new_n926), .A3(new_n938), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n793), .A2(new_n814), .ZN(new_n950));
  OAI21_X1  g525(.A(G290), .B1(new_n580), .B2(new_n584), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT104), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G303), .B(G305), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n956), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n954), .B1(new_n950), .B2(new_n951), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n942), .A2(new_n949), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n960), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT42), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(G868), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n963), .A2(KEYINPUT106), .A3(G868), .A4(new_n966), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n838), .A2(G868), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AND4_X1   g547(.A1(new_n918), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n967), .B2(new_n968), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n918), .B1(new_n974), .B2(new_n970), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n970), .ZN(G331));
  NAND2_X1  g552(.A1(G301), .A2(KEYINPUT108), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n979));
  NAND2_X1  g554(.A1(G171), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n538), .A2(new_n540), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n978), .B(new_n980), .C1(new_n530), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(G168), .A2(new_n979), .A3(G171), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n842), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n924), .A3(new_n983), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n938), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n943), .A3(new_n986), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n990), .B2(new_n964), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n961), .A3(new_n989), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n997));
  OR3_X1    g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n870), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT45), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n874), .B2(new_n861), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n1011));
  OR3_X1    g586(.A1(new_n1010), .A2(new_n1011), .A3(G1996), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1010), .B2(G1996), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n759), .B(G2067), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(new_n888), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1012), .B(new_n1013), .C1(new_n1010), .C2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n784), .A2(G1996), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1014), .B(new_n1020), .C1(new_n860), .C2(G1996), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1009), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT110), .Z(new_n1023));
  XOR2_X1   g598(.A(new_n801), .B(new_n804), .Z(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1009), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1010), .A2(G1986), .A3(G290), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT48), .Z(new_n1027));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n804), .ZN(new_n1028));
  OAI22_X1  g603(.A1(new_n1023), .A2(new_n1028), .B1(G2067), .B2(new_n875), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1025), .A2(new_n1027), .B1(new_n1029), .B2(new_n1009), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1018), .A2(new_n1019), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G290), .B(G1986), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1009), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1001), .B1(new_n494), .B2(new_n498), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1384), .B1(new_n861), .B2(new_n493), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT111), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G2084), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n870), .A2(new_n1041), .A3(new_n1001), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n870), .B2(new_n1001), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1040), .A2(KEYINPUT45), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n715), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1036), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT51), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1047), .A2(G168), .A3(new_n1051), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1054), .A2(new_n1056), .B1(G286), .B2(new_n1052), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(G8), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(KEYINPUT51), .C1(new_n1053), .C2(new_n1052), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT62), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(G286), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1036), .B1(new_n1005), .B2(new_n1045), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n814), .A2(G1976), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT114), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1071), .A3(new_n1068), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(KEYINPUT52), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n582), .A2(new_n1074), .A3(new_n585), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(KEYINPUT115), .A3(new_n1076), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  INV_X1    g658(.A(G1981), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n588), .A2(new_n1084), .A3(new_n592), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n588), .B2(new_n592), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1087), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT49), .A3(new_n1085), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1090), .A3(new_n1067), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1073), .A2(new_n1082), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1036), .B1(new_n514), .B2(new_n518), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n1094));
  OR3_X1    g669(.A1(new_n1093), .A2(new_n1094), .A3(KEYINPUT55), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(KEYINPUT55), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1093), .B2(KEYINPUT55), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1041), .B1(new_n870), .B2(new_n1001), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1045), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(G2090), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1040), .A2(KEYINPUT45), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1045), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n811), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1099), .B1(new_n1106), .B2(new_n1036), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1008), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1108));
  INV_X1    g683(.A(G2090), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1046), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n811), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1036), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1112), .A2(KEYINPUT113), .A3(new_n1098), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT113), .B1(new_n1112), .B2(new_n1098), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1092), .B(new_n1107), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1105), .B2(G2078), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1108), .A2(new_n1046), .ZN(new_n1119));
  INV_X1    g694(.A(G1961), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1045), .B(new_n1049), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(G2078), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(new_n1126), .A3(KEYINPUT123), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1961), .B1(new_n1108), .B2(new_n1046), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1118), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(G301), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1115), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1052), .A2(G168), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1115), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1112), .A2(new_n1098), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1138), .A2(new_n1136), .A3(new_n1135), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1139), .B(new_n1092), .C1(new_n1114), .C2(new_n1113), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1066), .A2(new_n1134), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1092), .ZN(new_n1143));
  AOI211_X1 g718(.A(G1976), .B(G288), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1067), .B1(new_n1144), .B2(new_n1086), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n545), .A2(KEYINPUT54), .A3(new_n549), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT54), .B1(new_n545), .B2(new_n549), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1103), .A2(new_n1045), .A3(new_n1124), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1007), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1121), .A2(KEYINPUT125), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1129), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .A4(new_n1117), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1149), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1132), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1064), .A2(new_n1115), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1956), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT56), .B(G2072), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1103), .A2(new_n1104), .A3(new_n1045), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT117), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT116), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1167), .A2(KEYINPUT116), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1168), .B(new_n1169), .C1(new_n929), .C2(new_n930), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n568), .A2(new_n572), .A3(KEYINPUT116), .A4(new_n1167), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1164), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(G1348), .B1(new_n1108), .B2(new_n1046), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n870), .A2(new_n1045), .A3(new_n1001), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(G2067), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1173), .B1(new_n612), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1160), .A2(new_n1162), .A3(new_n1171), .A4(new_n1170), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(G1341), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1175), .A2(KEYINPUT119), .A3(new_n1182), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1185), .B(new_n1186), .C1(G1996), .C2(new_n1105), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n557), .B1(new_n1188), .B2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT120), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1187), .A2(KEYINPUT120), .A3(new_n1191), .A4(new_n558), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1173), .A2(KEYINPUT61), .A3(new_n1179), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1177), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n612), .B1(new_n1177), .B2(KEYINPUT60), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT60), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1163), .A2(new_n1172), .ZN(new_n1203));
  AOI21_X1  g778(.A(KEYINPUT61), .B1(new_n1203), .B2(new_n1179), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT121), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1180), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1146), .B1(new_n1158), .B2(new_n1206), .ZN(new_n1207));
  AOI211_X1 g782(.A(new_n1032), .B(new_n1035), .C1(new_n1141), .C2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1158), .A2(new_n1206), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1146), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1057), .A2(KEYINPUT62), .A3(new_n1059), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1134), .B1(new_n1211), .B2(new_n1060), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1035), .ZN(new_n1215));
  AOI21_X1  g790(.A(KEYINPUT126), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1031), .B1(new_n1208), .B2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g792(.A1(G227), .A2(new_n460), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n1219), .B1(new_n660), .B2(new_n661), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1220), .B1(new_n703), .B2(new_n705), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1221), .B1(new_n995), .B2(new_n997), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n912), .B2(new_n914), .ZN(G308));
  NAND2_X1  g797(.A1(new_n912), .A2(new_n914), .ZN(new_n1224));
  OAI211_X1 g798(.A(new_n1224), .B(new_n1221), .C1(new_n997), .C2(new_n995), .ZN(G225));
endmodule


