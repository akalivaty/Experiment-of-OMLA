//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1187, new_n1188, new_n1189,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G107), .ZN(new_n232));
  INV_X1    g0032(.A(G264), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n213), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  OAI221_X1 g0035(.A(new_n216), .B1(new_n220), .B2(new_n223), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n235), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(new_n212), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n217), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n211), .B1(new_n206), .B2(new_n221), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n256), .A2(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n254), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n211), .A3(G1), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n218), .B1(new_n212), .B2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n267), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n210), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n264), .B1(G50), .B2(new_n267), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT9), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n218), .B1(new_n257), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n275), .A2(G274), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G226), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n279), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G223), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n284), .B1(new_n230), .B2(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n278), .B(new_n281), .C1(new_n287), .C2(new_n279), .ZN(new_n288));
  INV_X1    g0088(.A(G200), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n290), .A2(KEYINPUT66), .B1(G190), .B2(new_n288), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n273), .B(new_n291), .C1(KEYINPUT66), .C2(new_n290), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n272), .C1(G169), .C2(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT16), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT7), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G20), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n257), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT69), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT69), .A2(G33), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT73), .B(new_n303), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(KEYINPUT69), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT69), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT73), .B1(new_n312), .B2(new_n303), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n300), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT72), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n303), .A2(G33), .ZN(new_n317));
  AOI21_X1  g0117(.A(G20), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n318), .B2(KEYINPUT7), .ZN(new_n319));
  OAI211_X1 g0119(.A(KEYINPUT72), .B(new_n299), .C1(new_n282), .C2(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n202), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G58), .A2(G68), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n203), .A2(new_n205), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n261), .A2(G159), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(KEYINPUT71), .A3(G20), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n298), .B1(new_n322), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n310), .A2(KEYINPUT3), .A3(new_n311), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(new_n299), .A3(new_n211), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n211), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n202), .B1(new_n339), .B2(KEYINPUT7), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n330), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n268), .B1(new_n341), .B2(KEYINPUT16), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT74), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n298), .C1(new_n322), .C2(new_n330), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n332), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n256), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n270), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n269), .A2(new_n347), .B1(new_n267), .B2(new_n346), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(KEYINPUT75), .A3(new_n349), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n279), .A2(new_n277), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n278), .B1(G232), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G87), .ZN(new_n356));
  XOR2_X1   g0156(.A(new_n356), .B(KEYINPUT76), .Z(new_n357));
  NAND2_X1  g0157(.A1(new_n280), .A2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G223), .B2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n337), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n279), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G169), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n294), .B2(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n352), .A2(new_n353), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT18), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT78), .B1(new_n362), .B2(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n362), .A2(new_n289), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n355), .A2(new_n361), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n345), .A2(KEYINPUT79), .A3(new_n349), .A4(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT17), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n352), .A2(new_n377), .A3(new_n353), .A4(new_n366), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n368), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n259), .B2(new_n230), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n254), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT11), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n383), .A2(KEYINPUT67), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(KEYINPUT67), .ZN(new_n385));
  OR3_X1    g0185(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT12), .B1(new_n267), .B2(G68), .ZN(new_n387));
  INV_X1    g0187(.A(new_n269), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n202), .B1(new_n210), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n386), .A2(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n278), .B1(G238), .B2(new_n354), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n282), .A2(G232), .A3(G1698), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n282), .A2(G226), .A3(new_n283), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G97), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n275), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT13), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(KEYINPUT68), .A2(KEYINPUT14), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(G169), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n401), .B1(new_n398), .B2(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n391), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(G190), .ZN(new_n406));
  INV_X1    g0206(.A(new_n391), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n398), .A2(G200), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n346), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT15), .B(G87), .Z(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n259), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n254), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n270), .A2(G77), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(G77), .B2(new_n267), .C1(new_n269), .C2(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n279), .A2(new_n277), .A3(new_n231), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n232), .B2(new_n282), .C1(new_n285), .C2(new_n225), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n278), .B(new_n418), .C1(new_n420), .C2(new_n279), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n417), .B1(G190), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n289), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n294), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n417), .B(new_n424), .C1(G169), .C2(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n297), .A2(new_n379), .A3(new_n410), .A4(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n267), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n268), .B(new_n267), .C1(G1), .C2(new_n257), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n431), .B2(new_n428), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT81), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n314), .A2(new_n321), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n434), .A2(KEYINPUT80), .A3(new_n232), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT80), .B1(new_n434), .B2(new_n232), .ZN(new_n436));
  XOR2_X1   g0236(.A(G97), .B(G107), .Z(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT6), .A2(G97), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n437), .A2(KEYINPUT6), .B1(G107), .B2(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n433), .B1(new_n441), .B2(new_n254), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n275), .A2(G274), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n276), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n279), .B1(new_n446), .B2(new_n445), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G257), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n443), .A3(new_n451), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n455), .B(new_n456), .C1(new_n227), .C2(new_n285), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n333), .A2(new_n336), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G244), .A3(new_n283), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT4), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n453), .B(new_n454), .C1(new_n461), .C2(new_n275), .ZN(new_n462));
  INV_X1    g0262(.A(G169), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G179), .B2(new_n462), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n442), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n462), .A2(new_n372), .ZN(new_n467));
  INV_X1    g0267(.A(new_n454), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n452), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n461), .A2(new_n275), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n289), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n442), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n337), .A2(new_n475), .A3(G20), .A4(new_n226), .ZN(new_n476));
  INV_X1    g0276(.A(new_n282), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n211), .A2(G87), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n310), .B2(new_n311), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n211), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n232), .A2(KEYINPUT23), .A3(G20), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(new_n211), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n474), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n458), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n488));
  INV_X1    g0288(.A(new_n474), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n479), .A4(new_n485), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n268), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT25), .B1(new_n266), .B2(new_n232), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n232), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n430), .A2(new_n232), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n227), .A2(new_n283), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n458), .B(new_n496), .C1(G257), .C2(new_n283), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n312), .A2(G294), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n275), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n450), .A2(G264), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n499), .A2(new_n448), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G190), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n495), .B(new_n503), .C1(new_n289), .C2(new_n502), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n466), .A2(new_n473), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n431), .A2(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n266), .A2(new_n480), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n211), .A2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n254), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT85), .B1(new_n268), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n456), .B(new_n211), .C1(G33), .C2(new_n428), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n516), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n509), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G257), .A2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n233), .B2(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n458), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n477), .A2(G303), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n275), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n450), .A2(G270), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n449), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G169), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n506), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n526), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n448), .B1(G270), .B2(new_n450), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n534), .B(new_n521), .C1(new_n372), .C2(new_n533), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n519), .A2(new_n520), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n507), .A2(new_n508), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n529), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(KEYINPUT21), .A3(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n526), .A2(new_n528), .A3(new_n294), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AND4_X1   g0342(.A1(new_n530), .A2(new_n535), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n481), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n231), .A2(G1698), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G238), .B2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n337), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT84), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n279), .ZN(new_n549));
  INV_X1    g0349(.A(new_n446), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n275), .A2(G250), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n551), .B(KEYINPUT83), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n275), .A2(G274), .A3(new_n446), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n463), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n554), .B1(new_n548), .B2(new_n279), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n294), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n458), .A2(new_n211), .A3(G68), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n258), .A2(new_n561), .A3(G97), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n226), .B1(new_n395), .B2(new_n211), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n564), .B2(new_n561), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n268), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n266), .B2(new_n413), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n413), .B2(new_n430), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n557), .A2(new_n559), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n431), .A2(G87), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(G190), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n289), .C2(new_n558), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n497), .A2(new_n498), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n279), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(new_n294), .A3(new_n449), .A4(new_n500), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n502), .B2(G169), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n495), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n543), .A2(new_n569), .A3(new_n573), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n505), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n427), .A2(new_n581), .ZN(G372));
  AND3_X1   g0382(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n405), .B1(new_n583), .B2(new_n425), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n584), .A2(new_n376), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n350), .A2(new_n364), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n586), .B(new_n377), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n293), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n296), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n569), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT87), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT87), .B1(new_n569), .B2(new_n573), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n540), .A2(new_n530), .A3(new_n542), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n578), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n466), .A2(new_n473), .A3(new_n504), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n569), .A2(new_n573), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n442), .A2(new_n465), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n593), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT26), .B1(new_n466), .B2(new_n601), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n427), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n591), .A2(new_n609), .ZN(G369));
  NAND3_X1  g0410(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n611), .A2(KEYINPUT27), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(KEYINPUT27), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(G213), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(G343), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n521), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n596), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n535), .A2(new_n540), .A3(new_n530), .A4(new_n542), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n618), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G330), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n578), .A2(new_n617), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n616), .B1(new_n491), .B2(new_n494), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT88), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n628), .A2(new_n504), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n626), .B1(new_n630), .B2(new_n578), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n596), .A2(new_n617), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n626), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0439(.A(new_n214), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G41), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n563), .A2(new_n226), .A3(new_n480), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(G1), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n223), .B2(new_n642), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT28), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n499), .A2(new_n501), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n469), .A2(new_n470), .A3(new_n648), .A4(new_n541), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT90), .B1(new_n649), .B2(new_n556), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT30), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT30), .ZN(new_n652));
  OAI211_X1 g0452(.A(KEYINPUT90), .B(new_n652), .C1(new_n649), .C2(new_n556), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n449), .ZN(new_n654));
  AOI21_X1  g0454(.A(G179), .B1(new_n531), .B2(new_n532), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(new_n462), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n556), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n616), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT31), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(KEYINPUT31), .A3(new_n616), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(KEYINPUT91), .B1(new_n581), .B2(new_n617), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n665), .A3(new_n662), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n623), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT29), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n596), .A2(new_n578), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n603), .A3(new_n593), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n569), .B1(new_n670), .B2(new_n505), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n606), .A2(new_n607), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n668), .B(new_n617), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NOR4_X1   g0473(.A1(new_n601), .A2(new_n442), .A3(KEYINPUT26), .A4(new_n465), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n603), .A2(new_n605), .A3(new_n593), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n616), .B1(new_n600), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n673), .B1(new_n677), .B2(new_n668), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n647), .B1(new_n679), .B2(G1), .ZN(G364));
  XOR2_X1   g0480(.A(new_n624), .B(KEYINPUT92), .Z(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n265), .A2(G20), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n210), .B1(new_n683), .B2(G45), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n641), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n682), .B(new_n687), .C1(G330), .C2(new_n621), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n217), .B1(G20), .B2(new_n463), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT93), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n211), .A2(new_n294), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(G190), .A3(new_n289), .ZN(new_n695));
  INV_X1    g0495(.A(G322), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G190), .A2(G200), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G311), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n695), .A2(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n211), .A2(G179), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n697), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI211_X1 g0503(.A(new_n282), .B(new_n700), .C1(G329), .C2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(G190), .A3(G200), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G303), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n372), .A2(G179), .A3(G200), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n211), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n694), .A2(G200), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n372), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT94), .B(G326), .Z(new_n713));
  AOI22_X1  g0513(.A1(G294), .A2(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n711), .A2(G190), .ZN(new_n715));
  XNOR2_X1  g0515(.A(KEYINPUT33), .B(G317), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n701), .A2(new_n372), .A3(G200), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n715), .A2(new_n716), .B1(new_n718), .B2(G283), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n704), .A2(new_n707), .A3(new_n714), .A4(new_n719), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n226), .A2(new_n705), .B1(new_n717), .B2(new_n232), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(G50), .B2(new_n712), .ZN(new_n722));
  INV_X1    g0522(.A(G159), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n702), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT32), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n282), .B1(new_n695), .B2(new_n201), .ZN(new_n726));
  INV_X1    g0526(.A(new_n698), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n726), .B1(G77), .B2(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(G97), .A2(new_n710), .B1(new_n715), .B2(G68), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n722), .A2(new_n725), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n693), .B1(new_n720), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n214), .A2(new_n282), .ZN(new_n732));
  INV_X1    g0532(.A(G355), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(G116), .B2(new_n214), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n248), .A2(new_n276), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n337), .A2(new_n214), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n276), .B2(new_n222), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n692), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n686), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n741), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n621), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n688), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(G396));
  NAND2_X1  g0549(.A1(new_n693), .A2(new_n740), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n686), .B1(new_n750), .B2(G77), .ZN(new_n751));
  INV_X1    g0551(.A(G294), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n695), .A2(new_n752), .B1(new_n702), .B2(new_n699), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n282), .B(new_n753), .C1(G116), .C2(new_n727), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n706), .A2(G107), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G97), .A2(new_n710), .B1(new_n712), .B2(G303), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n715), .A2(G283), .B1(new_n718), .B2(G87), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n695), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G143), .B1(new_n727), .B2(G159), .ZN(new_n760));
  INV_X1    g0560(.A(new_n712), .ZN(new_n761));
  INV_X1    g0561(.A(G137), .ZN(new_n762));
  INV_X1    g0562(.A(new_n715), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n760), .B1(new_n761), .B2(new_n762), .C1(new_n260), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT34), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n706), .A2(G50), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n709), .A2(new_n201), .B1(new_n717), .B2(new_n202), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n337), .B(new_n768), .C1(G132), .C2(new_n703), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n764), .A2(new_n765), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n758), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n751), .B1(new_n772), .B2(new_n692), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n417), .A2(new_n616), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n423), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n425), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n425), .A2(new_n616), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n773), .B1(new_n779), .B2(new_n740), .ZN(new_n780));
  INV_X1    g0580(.A(new_n608), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n778), .B1(new_n781), .B2(new_n616), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n617), .B(new_n779), .C1(new_n671), .C2(new_n672), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n782), .A2(new_n667), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(new_n687), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n782), .A2(new_n783), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n667), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n780), .B1(new_n787), .B2(new_n790), .ZN(G384));
  AOI211_X1 g0591(.A(new_n480), .B(new_n220), .C1(new_n439), .C2(KEYINPUT35), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(KEYINPUT35), .B2(new_n439), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT36), .Z(new_n794));
  NAND3_X1  g0594(.A1(new_n222), .A2(G77), .A3(new_n323), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n221), .A2(G68), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n210), .B(G13), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n341), .A2(KEYINPUT16), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n348), .B1(new_n799), .B2(new_n342), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n614), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n801), .A2(KEYINPUT98), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT98), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n800), .B2(new_n614), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n379), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n352), .A2(new_n353), .A3(new_n802), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT37), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n345), .A2(new_n349), .A3(new_n374), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n367), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n801), .A2(new_n364), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n810), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT37), .B1(new_n806), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g0615(.A1(new_n807), .A2(KEYINPUT38), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT38), .B1(new_n807), .B2(new_n815), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT39), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n807), .A2(KEYINPUT38), .A3(new_n815), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n807), .A2(KEYINPUT101), .A3(KEYINPUT38), .A4(new_n815), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n808), .A2(new_n810), .A3(new_n586), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT37), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n825), .A2(new_n826), .A3(new_n811), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n825), .B2(new_n811), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n808), .B1(new_n587), .B2(new_n376), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n822), .B(new_n823), .C1(new_n830), .C2(KEYINPUT38), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n819), .B1(new_n831), .B2(new_n818), .ZN(new_n832));
  INV_X1    g0632(.A(new_n404), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n833), .A2(new_n400), .A3(new_n402), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n834), .A2(new_n391), .A3(new_n617), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT99), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n816), .A2(new_n817), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n391), .B(new_n616), .C1(new_n583), .C2(new_n834), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n391), .A2(new_n616), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n405), .A2(new_n409), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n783), .B2(new_n777), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT97), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n848), .A2(new_n849), .B1(new_n588), .B2(new_n614), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n838), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n590), .B1(new_n678), .B2(new_n427), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n851), .B(new_n852), .Z(new_n853));
  NAND2_X1  g0653(.A1(new_n662), .A2(KEYINPUT102), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n442), .A2(new_n472), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n605), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n601), .A2(new_n620), .A3(new_n578), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n504), .A4(new_n617), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n658), .A2(new_n859), .A3(KEYINPUT31), .A4(new_n616), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n854), .A2(new_n858), .A3(new_n661), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n778), .B1(new_n840), .B2(new_n842), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n822), .A2(new_n823), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n825), .A2(new_n811), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n829), .B1(new_n867), .B2(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n825), .A2(new_n826), .A3(new_n811), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n865), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n807), .A2(new_n815), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n863), .B1(new_n874), .B2(new_n820), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(KEYINPUT40), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n427), .A2(new_n861), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(G330), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n853), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n210), .B2(new_n683), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n853), .A2(new_n880), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n798), .B1(new_n882), .B2(new_n883), .ZN(G367));
  XOR2_X1   g0684(.A(new_n641), .B(KEYINPUT41), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n605), .A2(new_n616), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT104), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n856), .B1(new_n442), .B2(new_n617), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n637), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT44), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n637), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n893));
  XNOR2_X1  g0693(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n632), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT106), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n631), .B(new_n634), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n625), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n682), .B2(new_n899), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n679), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n891), .A2(new_n633), .A3(new_n894), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n895), .A2(KEYINPUT106), .A3(new_n632), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n898), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n885), .B1(new_n905), .B2(new_n679), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n685), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n889), .A2(new_n635), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n889), .A2(new_n578), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n616), .B1(new_n910), .B2(new_n466), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT43), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n571), .A2(new_n617), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n569), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT103), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n603), .A2(new_n593), .A3(new_n913), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n909), .A2(new_n911), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n912), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n919), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n889), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n633), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n907), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n244), .A2(new_n736), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n743), .B1(new_n640), .B2(new_n412), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n282), .B1(new_n717), .B2(new_n230), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT109), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n698), .A2(new_n221), .B1(new_n702), .B2(new_n762), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G150), .B2(new_n759), .ZN(new_n932));
  AOI22_X1  g0732(.A1(G143), .A2(new_n712), .B1(new_n715), .B2(G159), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n709), .A2(new_n202), .ZN(new_n934));
  INV_X1    g0734(.A(new_n705), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(G58), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n930), .A2(new_n932), .A3(new_n933), .A4(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n710), .A2(G107), .B1(new_n727), .B2(G283), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n761), .A2(new_n699), .B1(new_n717), .B2(new_n428), .ZN(new_n940));
  INV_X1    g0740(.A(G303), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n695), .A2(new_n941), .B1(new_n702), .B2(new_n942), .ZN(new_n943));
  NOR4_X1   g0743(.A1(new_n939), .A2(new_n940), .A3(new_n458), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n706), .A2(KEYINPUT46), .A3(G116), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n705), .A2(new_n480), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n945), .B1(KEYINPUT46), .B2(new_n946), .C1(new_n752), .C2(new_n763), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n944), .B1(KEYINPUT107), .B2(new_n938), .C1(new_n947), .C2(KEYINPUT108), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n937), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT47), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n692), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n686), .B1(new_n926), .B2(new_n928), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n918), .B2(new_n741), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n925), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(G387));
  NAND2_X1  g0757(.A1(new_n901), .A2(new_n685), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT110), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n901), .A2(new_n679), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n902), .A2(new_n960), .A3(new_n642), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n732), .A2(new_n644), .B1(G107), .B2(new_n214), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n241), .A2(new_n276), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n256), .A2(G50), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT50), .ZN(new_n965));
  AOI211_X1 g0765(.A(G45), .B(new_n643), .C1(G68), .C2(G77), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n736), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n962), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n686), .B1(new_n968), .B2(new_n743), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n705), .A2(new_n230), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G97), .B2(new_n718), .ZN(new_n971));
  XNOR2_X1  g0771(.A(KEYINPUT111), .B(G150), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n458), .C1(new_n702), .C2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT112), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n715), .A2(new_n346), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n759), .A2(G50), .B1(new_n727), .B2(G68), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n412), .A2(new_n710), .B1(new_n712), .B2(G159), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n458), .B1(new_n703), .B2(new_n713), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n759), .A2(G317), .B1(new_n727), .B2(G303), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n761), .B2(new_n696), .C1(new_n699), .C2(new_n763), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT48), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n710), .A2(G283), .B1(new_n935), .B2(G294), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT49), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n979), .B1(new_n480), .B2(new_n717), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n986), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(KEYINPUT49), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n978), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n969), .B1(new_n991), .B2(new_n692), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT113), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n631), .B2(new_n741), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n959), .A2(new_n961), .A3(new_n994), .ZN(G393));
  AND2_X1   g0795(.A1(new_n896), .A2(new_n903), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n905), .B(new_n641), .C1(new_n902), .C2(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n742), .B1(new_n428), .B2(new_n214), .C1(new_n251), .C2(new_n736), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n687), .B1(new_n998), .B2(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n703), .A2(G143), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n458), .B(new_n1000), .C1(new_n256), .C2(new_n698), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n763), .A2(new_n221), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n202), .A2(new_n705), .B1(new_n717), .B2(new_n226), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n709), .A2(new_n230), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n761), .A2(new_n260), .B1(new_n723), .B2(new_n695), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT51), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n761), .A2(new_n942), .B1(new_n699), .B2(new_n695), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT52), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n763), .A2(new_n941), .B1(new_n480), .B2(new_n709), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n477), .B1(new_n702), .B2(new_n696), .C1(new_n752), .C2(new_n698), .ZN(new_n1011));
  INV_X1    g0811(.A(G283), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n232), .A2(new_n717), .B1(new_n705), .B2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1005), .A2(new_n1007), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n999), .B1(KEYINPUT114), .B2(new_n998), .C1(new_n1015), .C2(new_n693), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n922), .B2(new_n741), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n996), .B2(new_n685), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n997), .A2(new_n1018), .ZN(G390));
  NAND2_X1  g0819(.A1(new_n861), .A2(G330), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n843), .A2(new_n779), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT115), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT115), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n861), .A2(new_n1023), .A3(G330), .A4(new_n862), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n845), .A2(new_n837), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n818), .B1(new_n866), .B2(new_n870), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n819), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n866), .A2(new_n870), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n777), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n677), .B2(new_n776), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n836), .B1(new_n1032), .B2(new_n844), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1025), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n650), .A2(KEYINPUT30), .B1(new_n656), .B2(new_n556), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n660), .B(new_n617), .C1(new_n1036), .C2(new_n653), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT31), .B1(new_n658), .B2(new_n616), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT91), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n666), .A2(new_n1039), .A3(new_n858), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1040), .A2(G330), .A3(new_n779), .A4(new_n843), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n836), .B1(new_n1032), .B2(new_n844), .C1(new_n866), .C2(new_n870), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n832), .C2(new_n1026), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1035), .A2(new_n685), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT117), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n427), .A2(G330), .A3(new_n861), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n852), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n783), .A2(new_n777), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n843), .B1(new_n667), .B2(new_n779), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n1025), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n779), .B1(new_n1020), .B2(KEYINPUT116), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT116), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n861), .B2(G330), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n844), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1041), .A2(new_n1032), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1048), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1046), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1035), .A2(new_n1043), .A3(new_n1058), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n641), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n686), .B1(new_n750), .B2(new_n346), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n695), .A2(new_n480), .B1(new_n702), .B2(new_n752), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n282), .B(new_n1064), .C1(G97), .C2(new_n727), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n706), .A2(G87), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1004), .B1(G68), .B2(new_n718), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G107), .A2(new_n715), .B1(new_n712), .B2(G283), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  INV_X1    g0870(.A(G125), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n698), .A2(new_n1070), .B1(new_n702), .B2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n477), .B(new_n1072), .C1(G132), .C2(new_n759), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n715), .A2(G137), .B1(new_n718), .B2(G50), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G159), .A2(new_n710), .B1(new_n712), .B2(G128), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n705), .A2(new_n972), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT53), .Z(new_n1078));
  OAI21_X1  g0878(.A(new_n1069), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1063), .B1(new_n1079), .B2(new_n692), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n832), .B2(new_n740), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n1045), .A2(new_n1062), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(G378));
  INV_X1    g0883(.A(new_n851), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n617), .B1(new_n1036), .B2(new_n653), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n859), .B1(new_n1085), .B2(KEYINPUT31), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n860), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1038), .B1(new_n581), .B2(new_n617), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1021), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n816), .B2(new_n817), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n623), .B1(new_n1091), .B2(new_n864), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT120), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1092), .A2(new_n871), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1092), .B2(new_n871), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n272), .A2(new_n802), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT119), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n297), .B(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1099));
  XOR2_X1   g0899(.A(new_n1098), .B(new_n1099), .Z(new_n1100));
  NOR3_X1   g0900(.A1(new_n1094), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1092), .A2(new_n871), .A3(new_n1093), .A4(new_n1100), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1084), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT121), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1090), .A2(KEYINPUT40), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n822), .A2(new_n823), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n868), .A2(new_n869), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n873), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1106), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(G330), .B1(new_n875), .B2(KEYINPUT40), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT120), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1092), .A2(new_n871), .A3(new_n1093), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1100), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n851), .A3(new_n1102), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1104), .A2(new_n1105), .A3(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1115), .A2(new_n851), .A3(KEYINPUT121), .A4(new_n1102), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n685), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1100), .A2(new_n739), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n686), .B1(new_n750), .B2(G50), .ZN(new_n1121));
  INV_X1    g0921(.A(G132), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n763), .A2(new_n1122), .B1(new_n761), .B2(new_n1071), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n759), .A2(G128), .B1(new_n727), .B2(G137), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n705), .B2(new_n1070), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(G150), .C2(new_n710), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n718), .A2(G159), .ZN(new_n1130));
  AOI211_X1 g0930(.A(G33), .B(G41), .C1(new_n703), .C2(G124), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n759), .A2(G107), .B1(new_n703), .B2(G283), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n413), .B2(new_n698), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1134), .A2(new_n934), .A3(new_n970), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n761), .A2(new_n480), .B1(new_n717), .B2(new_n201), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G97), .B2(new_n715), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n458), .A2(G41), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT58), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G50), .B(new_n1138), .C1(new_n257), .C2(new_n274), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT118), .Z(new_n1144));
  NAND4_X1  g0944(.A1(new_n1132), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1121), .B1(new_n1145), .B2(new_n692), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1120), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1119), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1048), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1061), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1117), .A2(new_n1150), .A3(new_n1118), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1115), .A2(new_n851), .A3(new_n1102), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n851), .B1(new_n1115), .B2(new_n1102), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1150), .B(KEYINPUT57), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n641), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(G375));
  NAND2_X1  g0959(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n844), .A2(new_n739), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n686), .B1(new_n750), .B2(G68), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n761), .A2(new_n1122), .B1(new_n221), .B2(new_n709), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n763), .A2(new_n1070), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n706), .A2(G159), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n698), .A2(new_n260), .B1(new_n702), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G137), .B2(new_n759), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n337), .B1(G58), .B2(new_n718), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1166), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n695), .A2(new_n1012), .B1(new_n702), .B2(new_n941), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n282), .B(new_n1172), .C1(G107), .C2(new_n727), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n706), .A2(G97), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n710), .A2(new_n412), .B1(new_n718), .B2(G77), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G116), .A2(new_n715), .B1(new_n712), .B2(G294), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1162), .B1(new_n1178), .B2(new_n692), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1160), .A2(new_n685), .B1(new_n1161), .B2(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1058), .A2(new_n885), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1160), .A2(new_n1149), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(G381));
  NOR4_X1   g0983(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n956), .A2(new_n1184), .ZN(new_n1185));
  OR4_X1    g0985(.A1(G378), .A2(G375), .A3(new_n1185), .A4(G381), .ZN(G407));
  NAND2_X1  g0986(.A1(new_n615), .A2(G213), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT122), .Z(new_n1188));
  NAND3_X1  g0988(.A1(new_n1158), .A2(new_n1082), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(G407), .A2(G213), .A3(new_n1189), .ZN(G409));
  OR2_X1    g0990(.A1(new_n1151), .A2(new_n885), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n685), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1192), .A2(new_n1147), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G378), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1158), .B2(G378), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1156), .A2(new_n641), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1152), .B2(new_n1151), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1199), .A2(KEYINPUT123), .A3(new_n1148), .A4(new_n1082), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1195), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1188), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1059), .A2(KEYINPUT60), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1059), .A2(new_n1182), .A3(KEYINPUT60), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n641), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1180), .ZN(new_n1207));
  INV_X1    g1007(.A(G384), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(G384), .A3(new_n1180), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1201), .A2(KEYINPUT62), .A3(new_n1202), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1148), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(G378), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT123), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1158), .A2(new_n1196), .A3(G378), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1194), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1187), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1212), .B1(new_n1221), .B2(KEYINPUT62), .ZN(new_n1222));
  INV_X1    g1022(.A(G2897), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1220), .A2(new_n1223), .A3(new_n1187), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1209), .A2(new_n1210), .B1(G2897), .B2(new_n1188), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT127), .B1(new_n1227), .B2(KEYINPUT61), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1218), .B2(new_n1188), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT127), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT61), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1222), .A2(new_n1228), .A3(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n907), .A2(new_n924), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT124), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n955), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G390), .A2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(G393), .B(new_n748), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n956), .C2(new_n1240), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G390), .B1(new_n956), .B2(KEYINPUT125), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1242), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n956), .A2(KEYINPUT125), .A3(G390), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1243), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1234), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1229), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1220), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1201), .A2(new_n1202), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1247), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1245), .A3(new_n1244), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1243), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1251), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1219), .B1(new_n1259), .B2(new_n1195), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT63), .B1(new_n1260), .B2(new_n1211), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT126), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1248), .A2(new_n1232), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1201), .A2(new_n1187), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1229), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1201), .A2(new_n1187), .A3(new_n1211), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1252), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .A4(new_n1254), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1250), .A2(new_n1270), .ZN(G405));
  OAI21_X1  g1071(.A(new_n1259), .B1(G378), .B2(new_n1158), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(new_n1211), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(new_n1249), .ZN(G402));
endmodule


