//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT87), .ZN(new_n209));
  OR2_X1    g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n203), .A2(new_n204), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n214), .B1(new_n212), .B2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n207), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n209), .A2(new_n213), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT15), .B(new_n212), .C1(new_n208), .C2(new_n214), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G15gat), .B(G22gat), .Z(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(KEYINPUT16), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n223), .A2(new_n226), .A3(KEYINPUT89), .A4(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n224), .A2(G1gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(new_n224), .B2(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(KEYINPUT88), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n227), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT90), .B(new_n220), .C1(new_n232), .C2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n232), .A2(new_n237), .ZN(new_n240));
  INV_X1    g039(.A(new_n220), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n220), .B1(new_n232), .B2(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n238), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(new_n218), .B2(new_n219), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n249), .A3(new_n219), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n240), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT18), .A3(new_n246), .A4(new_n243), .ZN(new_n255));
  INV_X1    g054(.A(new_n252), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  INV_X1    g056(.A(new_n240), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n246), .B(new_n243), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n248), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G141gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G169gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G197gat), .ZN(new_n268));
  INV_X1    g067(.A(G169gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n266), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G197gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n263), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n272), .A3(new_n263), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n276), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT86), .B1(new_n278), .B2(new_n273), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n276), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n248), .A2(new_n261), .A3(new_n255), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n286));
  INV_X1    g085(.A(G211gat), .ZN(new_n287));
  INV_X1    g086(.A(G218gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(KEYINPUT22), .B2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G211gat), .B(G218gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT3), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n298), .B2(KEYINPUT2), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(G141gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G148gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n295), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n294), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(KEYINPUT80), .ZN(new_n314));
  AND2_X1   g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n313), .B2(KEYINPUT80), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT75), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n292), .B1(new_n320), .B2(new_n293), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n294), .A2(new_n308), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n323), .B(KEYINPUT81), .Z(new_n324));
  OAI21_X1  g123(.A(new_n315), .B1(new_n324), .B2(new_n321), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G78gat), .B(G106gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT79), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT31), .B(G50gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G22gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n325), .A3(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n269), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n336), .B2(KEYINPUT23), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT65), .B(G183gat), .Z(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT24), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n344), .B2(new_n346), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n341), .B(new_n343), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT64), .B(G169gat), .Z(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT23), .A3(new_n338), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n355), .A3(new_n341), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n342), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT28), .A3(new_n346), .ZN(new_n360));
  NOR2_X1   g159(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT65), .B(G183gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(KEYINPUT27), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n364), .B2(KEYINPUT28), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n337), .B1(new_n339), .B2(KEYINPUT26), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(KEYINPUT26), .B2(new_n337), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n348), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(new_n293), .B1(G226gat), .B2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(G226gat), .A3(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n292), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n372), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n292), .B1(new_n375), .B2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G8gat), .B(G36gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT71), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(KEYINPUT30), .A3(new_n382), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n381), .B(KEYINPUT72), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G113gat), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n393), .A2(G120gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(G120gat), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT1), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G127gat), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n391), .A2(new_n397), .A3(G134gat), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n390), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(KEYINPUT3), .B2(new_n311), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT75), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(new_n308), .B2(new_n318), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n310), .A2(new_n401), .A3(new_n312), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n308), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT76), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(KEYINPUT5), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n406), .A2(new_n409), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n412), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n406), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n407), .B2(KEYINPUT4), .ZN(new_n418));
  INV_X1    g217(.A(new_n401), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n419), .A2(KEYINPUT4), .A3(new_n311), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n407), .A2(new_n417), .A3(KEYINPUT4), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n401), .B(new_n308), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n412), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n414), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT0), .ZN(new_n429));
  XNOR2_X1  g228(.A(G57gat), .B(G85gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT83), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n412), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n412), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT39), .B1(new_n424), .B2(new_n412), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n434), .B(new_n437), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n438), .B(KEYINPUT39), .C1(new_n412), .C2(new_n424), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n434), .A4(new_n437), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n389), .A2(new_n433), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n414), .B(new_n431), .C1(new_n423), .C2(new_n426), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n431), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n427), .A2(new_n453), .A3(KEYINPUT6), .A4(new_n450), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n377), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT37), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n381), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT38), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n387), .A2(KEYINPUT38), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n383), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n335), .B(new_n446), .C1(new_n455), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n335), .A2(KEYINPUT82), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n333), .A2(new_n466), .A3(new_n334), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n447), .ZN(new_n469));
  INV_X1    g268(.A(new_n422), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n470), .A2(new_n418), .A3(new_n420), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT5), .B(new_n425), .C1(new_n471), .C2(new_n416), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n431), .B1(new_n472), .B2(new_n414), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n451), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n389), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT68), .ZN(new_n479));
  XOR2_X1   g278(.A(G71gat), .B(G99gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n369), .A2(new_n401), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n358), .A2(new_n368), .A3(new_n419), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  INV_X1    g283(.A(G233gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT33), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n487), .B(KEYINPUT32), .C1(new_n488), .C2(new_n481), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n486), .B(new_n495), .C1(new_n482), .C2(new_n483), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n491), .A3(new_n492), .ZN(new_n502));
  NAND2_X1  g301(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n503), .B1(new_n501), .B2(new_n502), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n464), .A2(new_n477), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n335), .A2(new_n501), .A3(new_n502), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n385), .A2(new_n388), .A3(new_n513), .A4(new_n386), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n455), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n476), .B2(new_n512), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n285), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G57gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT92), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G57gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n523), .A3(G64gat), .ZN(new_n524));
  INV_X1    g323(.A(G64gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G57gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT92), .B(G57gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT93), .A3(G64gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(KEYINPUT91), .A3(new_n533), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n520), .A2(G64gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n531), .A2(new_n539), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n258), .B1(KEYINPUT21), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT94), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n544), .A2(KEYINPUT21), .ZN(new_n548));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G127gat), .B(G155gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  XOR2_X1   g354(.A(G183gat), .B(G211gat), .Z(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n547), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n546), .A3(new_n557), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n564), .A2(new_n567), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n563), .ZN(new_n573));
  NOR2_X1   g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT97), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576));
  INV_X1    g375(.A(G99gat), .ZN(new_n577));
  INV_X1    g376(.A(G106gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n579), .B2(new_n563), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n572), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n571), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT97), .B1(new_n573), .B2(new_n574), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n576), .A3(new_n563), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n220), .A2(new_n589), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n257), .B2(new_n589), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT96), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT95), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n560), .A2(new_n562), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n544), .A2(new_n589), .A3(KEYINPUT10), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n544), .A2(new_n589), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n544), .A2(new_n589), .A3(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n544), .B2(new_n589), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n581), .A2(new_n588), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n530), .B2(new_n528), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n543), .A2(new_n540), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT98), .B(new_n614), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n610), .A2(new_n611), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n620));
  AOI21_X1  g419(.A(new_n607), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n605), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n610), .A2(new_n611), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n613), .A2(new_n618), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n606), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(KEYINPUT101), .A3(new_n622), .ZN(new_n629));
  INV_X1    g428(.A(new_n619), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n623), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n624), .A2(new_n629), .A3(new_n631), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n623), .ZN(new_n637));
  INV_X1    g436(.A(new_n631), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n604), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n519), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n474), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n222), .ZN(G1324gat));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n475), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT42), .B1(new_n645), .B2(new_n227), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT16), .B(G8gat), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g447(.A(KEYINPUT42), .B(new_n646), .S(new_n648), .Z(G1325gat));
  INV_X1    g448(.A(new_n501), .ZN(new_n650));
  INV_X1    g449(.A(new_n502), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n642), .A2(G15gat), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  INV_X1    g454(.A(new_n509), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n507), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT102), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n519), .A2(new_n641), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n654), .B1(G15gat), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT103), .Z(G1326gat));
  INV_X1    g461(.A(new_n468), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n560), .A2(new_n562), .ZN(new_n667));
  INV_X1    g466(.A(new_n603), .ZN(new_n668));
  INV_X1    g467(.A(new_n640), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT104), .Z(new_n671));
  AND2_X1   g470(.A1(new_n671), .A2(new_n519), .ZN(new_n672));
  INV_X1    g471(.A(new_n474), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n203), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n511), .A2(new_n518), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n603), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n560), .A2(new_n562), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n560), .B2(new_n562), .ZN(new_n682));
  NOR4_X1   g481(.A1(new_n681), .A2(new_n682), .A3(new_n285), .A4(new_n640), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n464), .B(new_n477), .C1(new_n658), .C2(new_n657), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n603), .B1(new_n684), .B2(new_n518), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n679), .B(new_n683), .C1(new_n685), .C2(KEYINPUT44), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n474), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n675), .A2(new_n687), .ZN(G1328gat));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n204), .A3(new_n389), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(KEYINPUT46), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT106), .Z(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n686), .B2(new_n475), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(KEYINPUT46), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(G1329gat));
  INV_X1    g493(.A(G43gat), .ZN(new_n695));
  INV_X1    g494(.A(new_n659), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n686), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(G43gat), .B1(new_n672), .B2(new_n652), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT47), .Z(G1330gat));
  XOR2_X1   g499(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n701));
  OAI211_X1 g500(.A(KEYINPUT108), .B(G50gat), .C1(new_n686), .C2(new_n663), .ZN(new_n702));
  INV_X1    g501(.A(G50gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n672), .A2(new_n703), .A3(new_n468), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n335), .A2(new_n501), .A3(new_n502), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n474), .A3(new_n475), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n707), .A2(KEYINPUT35), .B1(new_n455), .B2(new_n515), .ZN(new_n708));
  INV_X1    g507(.A(new_n463), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n709), .A2(new_n454), .A3(new_n449), .A4(new_n452), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n446), .A2(new_n335), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n710), .A2(new_n711), .B1(new_n476), .B2(new_n468), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n708), .B1(new_n712), .B2(new_n696), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n677), .B1(new_n713), .B2(new_n603), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n714), .A2(new_n468), .A3(new_n679), .A4(new_n683), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT108), .B1(new_n715), .B2(G50gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n701), .B1(new_n705), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G50gat), .B1(new_n686), .B2(new_n335), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(KEYINPUT48), .A3(new_n704), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(KEYINPUT109), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(new_n713), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n604), .A2(new_n284), .A3(new_n669), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n474), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n529), .ZN(G1332gat));
  INV_X1    g528(.A(new_n727), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n475), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT110), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n732), .B(new_n734), .ZN(G1333gat));
  NAND3_X1  g534(.A1(new_n730), .A2(G71gat), .A3(new_n659), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n727), .A2(new_n653), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(G71gat), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n730), .A2(new_n468), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  INV_X1    g540(.A(new_n667), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n284), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n640), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT111), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n714), .A2(new_n679), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n474), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n685), .A2(new_n743), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n685), .A2(KEYINPUT51), .A3(new_n743), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n673), .A2(new_n568), .A3(new_n640), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT112), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n747), .B1(new_n752), .B2(new_n754), .ZN(G1336gat));
  AOI21_X1  g554(.A(new_n669), .B1(new_n750), .B2(new_n751), .ZN(new_n756));
  AOI21_X1  g555(.A(G92gat), .B1(new_n756), .B2(new_n389), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n746), .A2(new_n569), .A3(new_n475), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT52), .ZN(G1337gat));
  AOI21_X1  g559(.A(G99gat), .B1(new_n756), .B2(new_n652), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n577), .A3(new_n696), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT113), .ZN(G1338gat));
  NAND4_X1  g563(.A1(new_n756), .A2(new_n578), .A3(new_n334), .A4(new_n333), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT114), .B(G106gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n746), .B2(new_n335), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n746), .B2(new_n663), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(new_n768), .ZN(G1339gat));
  NOR3_X1   g571(.A1(new_n604), .A2(new_n284), .A3(new_n640), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n681), .A2(new_n682), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n621), .B2(new_n623), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n624), .A2(new_n776), .A3(new_n629), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n635), .B1(new_n637), .B2(new_n775), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT55), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n636), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n268), .A2(new_n272), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n245), .A2(new_n247), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n246), .B1(new_n254), .B2(new_n243), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n283), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT55), .B1(new_n777), .B2(new_n778), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n668), .A2(new_n780), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n640), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n779), .A2(new_n284), .A3(new_n636), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n787), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n792), .B2(new_n668), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n773), .B1(new_n774), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n794), .A2(new_n474), .A3(new_n389), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n706), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT115), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n284), .A2(new_n393), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT116), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n468), .A2(new_n653), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n285), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1340gat));
  INV_X1    g603(.A(G120gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n805), .A3(new_n640), .ZN(new_n806));
  OAI21_X1  g605(.A(G120gat), .B1(new_n802), .B2(new_n669), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT117), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1341gat));
  OAI21_X1  g611(.A(G127gat), .B1(new_n802), .B2(new_n774), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n742), .A2(new_n397), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n796), .B2(new_n814), .ZN(G1342gat));
  NOR2_X1   g614(.A1(new_n794), .A2(new_n474), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n389), .A2(new_n603), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n801), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G134gat), .ZN(new_n820));
  INV_X1    g619(.A(G134gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n821), .A3(new_n706), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n822), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT118), .B1(new_n822), .B2(KEYINPUT56), .ZN(new_n824));
  OAI221_X1 g623(.A(new_n820), .B1(KEYINPUT56), .B2(new_n822), .C1(new_n823), .C2(new_n824), .ZN(G1343gat));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n335), .B(new_n659), .C1(new_n816), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT120), .B1(new_n794), .B2(new_n474), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(new_n302), .A3(new_n475), .A4(new_n284), .ZN(new_n830));
  INV_X1    g629(.A(new_n300), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n794), .A2(KEYINPUT57), .A3(new_n335), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n696), .A2(new_n673), .A3(new_n475), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n777), .A2(KEYINPUT119), .A3(new_n778), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT119), .B1(new_n777), .B2(new_n778), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n790), .B1(new_n838), .B2(new_n791), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n788), .B1(new_n839), .B2(new_n668), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n773), .B1(new_n667), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n841), .B2(new_n663), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n831), .B1(new_n843), .B2(new_n285), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n830), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n847), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n669), .A2(G148gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n827), .A2(new_n475), .A3(new_n828), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT121), .Z(new_n852));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(G148gat), .C1(new_n843), .C2(new_n669), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT122), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n663), .A2(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT123), .B(new_n788), .C1(new_n839), .C2(new_n668), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n742), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n773), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n794), .B2(new_n335), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n833), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n640), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n853), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n852), .B1(new_n855), .B2(new_n866), .ZN(G1345gat));
  NAND4_X1  g666(.A1(new_n829), .A2(new_n296), .A3(new_n475), .A4(new_n742), .ZN(new_n868));
  OAI21_X1  g667(.A(G155gat), .B1(new_n843), .B2(new_n774), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  NAND3_X1  g669(.A1(new_n829), .A2(new_n297), .A3(new_n817), .ZN(new_n871));
  OAI21_X1  g670(.A(G162gat), .B1(new_n843), .B2(new_n603), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1347gat));
  NAND2_X1  g672(.A1(new_n474), .A2(new_n389), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n794), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n801), .ZN(new_n876));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876), .B2(new_n285), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n706), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n284), .A2(new_n354), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(G1348gat));
  OAI21_X1  g679(.A(G176gat), .B1(new_n876), .B2(new_n669), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n640), .A2(new_n338), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1349gat));
  OAI21_X1  g682(.A(new_n362), .B1(new_n876), .B2(new_n774), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n742), .A2(new_n359), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g686(.A1(new_n878), .A2(G190gat), .A3(new_n603), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT124), .ZN(new_n889));
  OAI21_X1  g688(.A(G190gat), .B1(new_n876), .B2(new_n603), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(G1351gat));
  NAND4_X1  g693(.A1(new_n875), .A2(new_n334), .A3(new_n333), .A4(new_n696), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n284), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n659), .A2(new_n874), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n863), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n285), .A2(new_n271), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n898), .A2(new_n271), .B1(new_n900), .B2(new_n901), .ZN(G1352gat));
  NOR3_X1   g701(.A1(new_n895), .A2(G204gat), .A3(new_n669), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT62), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n863), .A2(new_n640), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G204gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1353gat));
  NAND4_X1  g706(.A1(new_n861), .A2(new_n742), .A3(new_n862), .A4(new_n899), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(G211gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n896), .A2(new_n287), .A3(new_n742), .A4(new_n897), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT127), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1354gat));
  NAND4_X1  g721(.A1(new_n896), .A2(new_n288), .A3(new_n668), .A4(new_n897), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n900), .A2(new_n668), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n288), .ZN(G1355gat));
endmodule


