//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  OAI211_X1 g002(.A(new_n187), .B(G146), .C1(new_n188), .C2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT71), .A3(new_n191), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT68), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT68), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n201), .B1(new_n204), .B2(G137), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n200), .B1(new_n202), .B2(new_n203), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n205), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n200), .A2(G134), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n216), .B2(G131), .ZN(new_n217));
  AOI211_X1 g031(.A(KEYINPUT70), .B(new_n211), .C1(new_n206), .C2(new_n215), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n199), .B(new_n212), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT68), .A2(G134), .ZN(new_n225));
  AOI21_X1  g039(.A(G137), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n226), .B2(new_n214), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT70), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n213), .A3(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(KEYINPUT72), .A3(new_n199), .A4(new_n212), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n190), .A2(G143), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n187), .A2(G146), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n187), .A2(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n190), .A2(G143), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT66), .A3(KEYINPUT0), .A4(G128), .ZN(new_n240));
  OR3_X1    g054(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n236), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n225), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n245), .A2(new_n200), .B1(new_n207), .B2(new_n208), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n224), .A2(G137), .A3(new_n225), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT69), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n246), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n205), .B2(new_n210), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n221), .A2(new_n231), .A3(KEYINPUT30), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G116), .B(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n256), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n219), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n255), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n262), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n221), .A2(new_n231), .A3(new_n267), .A4(new_n254), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n251), .B1(new_n246), .B2(new_n249), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n205), .A2(new_n210), .A3(new_n250), .ZN(new_n279));
  INV_X1    g093(.A(new_n242), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n196), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n241), .B1(new_n234), .B2(new_n235), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n278), .A2(new_n279), .B1(new_n282), .B2(new_n240), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n217), .A2(new_n218), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n199), .A2(new_n212), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n286), .B2(KEYINPUT72), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n287), .A2(KEYINPUT28), .A3(new_n267), .A4(new_n221), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n267), .B1(new_n254), .B2(new_n219), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n254), .A2(new_n219), .A3(new_n267), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n274), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n276), .A2(new_n277), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n276), .A2(new_n296), .A3(new_n277), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n290), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n231), .A2(new_n254), .ZN(new_n300));
  INV_X1    g114(.A(new_n221), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n262), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n268), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n275), .A2(new_n277), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n295), .A2(new_n297), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n310), .B(new_n274), .C1(new_n288), .C2(new_n292), .ZN(new_n311));
  INV_X1    g125(.A(new_n289), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n298), .B(new_n312), .C1(new_n268), .C2(new_n290), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT74), .B1(new_n313), .B2(new_n275), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n266), .A2(new_n274), .A3(new_n268), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT31), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n266), .A2(new_n318), .A3(new_n274), .A4(new_n268), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n315), .B(new_n317), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G472), .A2(G902), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n309), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n319), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n313), .A2(new_n275), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n310), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n313), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n317), .A3(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n309), .B(new_n323), .C1(new_n326), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n308), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G237), .ZN(new_n334));
  INV_X1    g148(.A(G953), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G214), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n187), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n270), .A2(G143), .A3(G214), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT18), .A3(G131), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G125), .ZN(new_n342));
  INV_X1    g156(.A(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n190), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT18), .A2(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n337), .A2(new_n338), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n340), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G113), .B(G122), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT88), .B(G104), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n270), .A2(G143), .A3(G214), .ZN(new_n356));
  AOI21_X1  g170(.A(G143), .B1(new_n270), .B2(G214), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT17), .B(G131), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT89), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n339), .A2(new_n360), .A3(KEYINPUT17), .A4(G131), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT16), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n343), .A2(KEYINPUT16), .A3(G140), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT78), .A4(G146), .ZN(new_n365));
  AOI21_X1  g179(.A(G146), .B1(new_n363), .B2(new_n364), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n364), .A3(G146), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n362), .A2(KEYINPUT90), .A3(new_n365), .A4(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n339), .B(new_n211), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n363), .A2(new_n364), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n190), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n375), .A2(new_n365), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT90), .B1(new_n378), .B2(new_n362), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n351), .B(new_n355), .C1(new_n374), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n362), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n373), .A3(new_n370), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(KEYINPUT91), .A3(new_n351), .A4(new_n355), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n351), .B1(new_n374), .B2(new_n379), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT92), .B1(new_n389), .B2(new_n354), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(KEYINPUT92), .A3(new_n354), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G902), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  INV_X1    g210(.A(new_n371), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n345), .B1(KEYINPUT87), .B2(KEYINPUT19), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n399));
  MUX2_X1   g213(.A(new_n345), .B(new_n398), .S(new_n399), .Z(new_n400));
  OAI211_X1 g214(.A(new_n397), .B(new_n368), .C1(new_n400), .C2(G146), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n355), .B1(new_n401), .B2(new_n351), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n382), .B2(new_n387), .ZN(new_n408));
  INV_X1    g222(.A(new_n406), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT20), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G122), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G116), .ZN(new_n413));
  INV_X1    g227(.A(G116), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G122), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n187), .A2(G128), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT13), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n188), .A2(G143), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n419), .A2(new_n420), .ZN(new_n424));
  OAI21_X1  g238(.A(G134), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n204), .A2(new_n419), .A3(new_n422), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n417), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n419), .A2(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n245), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n432), .A2(new_n413), .A3(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n428), .B(new_n431), .C1(new_n434), .C2(new_n417), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT9), .B(G234), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(G953), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n427), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n427), .B2(new_n435), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n394), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT94), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n444), .A3(new_n394), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G478), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n448), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n396), .A2(new_n411), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n417), .A2(G104), .ZN(new_n454));
  AND2_X1   g268(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n455));
  NOR2_X1   g269(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G104), .B(G107), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n455), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G101), .ZN(new_n461));
  INV_X1    g275(.A(G101), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n457), .B(new_n462), .C1(new_n455), .C2(new_n458), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT4), .ZN(new_n464));
  XOR2_X1   g278(.A(G104), .B(G107), .Z(new_n465));
  INV_X1    g279(.A(new_n455), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n462), .B1(new_n467), .B2(new_n457), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n262), .B(new_n461), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(G101), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n414), .A2(KEYINPUT5), .A3(G119), .ZN(new_n473));
  INV_X1    g287(.A(G113), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n472), .A2(new_n475), .B1(new_n257), .B2(new_n258), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G122), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n469), .A2(new_n477), .A3(new_n479), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n478), .B(new_n480), .C1(KEYINPUT83), .C2(new_n483), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n244), .A2(G125), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n199), .A2(new_n343), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n335), .A2(G224), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n487), .A2(new_n488), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n463), .A2(new_n470), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n258), .A2(new_n497), .A3(KEYINPUT5), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n475), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n499), .B2(new_n259), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n479), .B(KEYINPUT8), .Z(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n476), .B2(new_n495), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n493), .A2(new_n494), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n494), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT85), .B1(new_n489), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n489), .A2(KEYINPUT85), .A3(new_n505), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n504), .B(new_n482), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n492), .A2(new_n394), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n492), .A2(new_n509), .A3(new_n394), .A4(new_n511), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT86), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n516), .A3(new_n512), .ZN(new_n517));
  NAND2_X1  g331(.A1(G234), .A2(G237), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(G952), .A3(new_n335), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(G902), .A3(G953), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G214), .B1(G237), .B2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n515), .A2(new_n517), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT10), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n192), .A2(new_n193), .B1(new_n197), .B2(new_n196), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(new_n195), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n198), .A2(new_n189), .A3(new_n191), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n463), .A3(new_n470), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n532), .A2(new_n471), .B1(new_n534), .B2(new_n530), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n244), .B(new_n461), .C1(new_n464), .C2(new_n468), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n535), .A2(new_n536), .B1(new_n278), .B2(new_n279), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n278), .A2(new_n279), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT82), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT82), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n278), .A2(new_n279), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n535), .A2(new_n536), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n335), .A2(G227), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT80), .ZN(new_n545));
  XNOR2_X1  g359(.A(G110), .B(G140), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n538), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n535), .A2(new_n536), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n540), .A2(new_n542), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n534), .B1(new_n471), .B2(new_n199), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n539), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n539), .A3(KEYINPUT12), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n550), .A2(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n548), .B(G469), .C1(new_n557), .C2(new_n547), .ZN(new_n558));
  INV_X1    g372(.A(G469), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(new_n394), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n547), .ZN(new_n563));
  INV_X1    g377(.A(new_n543), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n537), .ZN(new_n565));
  INV_X1    g379(.A(new_n556), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT12), .B1(new_n552), .B2(new_n539), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n543), .B(new_n547), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(G469), .B(G902), .C1(new_n565), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n529), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n453), .A2(new_n528), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n437), .B1(G234), .B2(new_n394), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n335), .A2(G221), .A3(G234), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  NAND2_X1  g390(.A1(new_n188), .A2(G119), .ZN(new_n577));
  INV_X1    g391(.A(G119), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G128), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT24), .B(G110), .ZN(new_n581));
  OR3_X1    g395(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT76), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT76), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n579), .A2(KEYINPUT23), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT77), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT23), .ZN(new_n587));
  OAI22_X1  g401(.A1(new_n584), .A2(new_n585), .B1(new_n587), .B2(new_n577), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n582), .A2(new_n583), .B1(new_n588), .B2(G110), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n375), .A2(new_n365), .A3(new_n377), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n580), .A2(new_n581), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n588), .B2(G110), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n368), .A3(new_n347), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT79), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n591), .B2(new_n594), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n576), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n576), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n595), .B2(KEYINPUT79), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n394), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT25), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n599), .A2(KEYINPUT25), .A3(new_n394), .A4(new_n601), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n573), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n599), .A2(new_n601), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(G902), .A3(new_n572), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n333), .A2(new_n571), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  OAI21_X1  g425(.A(KEYINPUT33), .B1(new_n440), .B2(KEYINPUT97), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n441), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G478), .ZN(new_n614));
  INV_X1    g428(.A(G478), .ZN(new_n615));
  MUX2_X1   g429(.A(new_n394), .B(new_n442), .S(new_n615), .Z(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n396), .B2(new_n411), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n513), .A2(new_n619), .A3(new_n514), .ZN(new_n620));
  INV_X1    g434(.A(new_n524), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n495), .A2(new_n476), .ZN(new_n622));
  INV_X1    g436(.A(new_n502), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n489), .A2(new_n505), .B1(new_n624), .B2(new_n500), .ZN(new_n625));
  INV_X1    g439(.A(new_n506), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n507), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n627), .B2(new_n482), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT96), .A3(new_n511), .A4(new_n492), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n620), .A2(new_n525), .A3(new_n621), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n618), .A2(new_n631), .A3(KEYINPUT98), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT98), .B1(new_n618), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n323), .B1(new_n326), .B2(new_n330), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n322), .B2(new_n394), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT95), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n394), .B1(new_n326), .B2(new_n330), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G472), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n609), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n634), .A2(new_n644), .A3(new_n645), .A4(new_n570), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT34), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n450), .A2(new_n451), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n396), .A2(new_n411), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n630), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n645), .A2(new_n570), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n640), .A2(new_n643), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n600), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n595), .B(new_n656), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n657), .A2(new_n394), .A3(new_n573), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n604), .A2(new_n605), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(new_n572), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n570), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n663), .A2(new_n453), .A3(new_n528), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n643), .A3(new_n640), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n635), .A2(KEYINPUT32), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n331), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n663), .B1(new_n669), .B2(new_n308), .ZN(new_n670));
  AOI22_X1  g484(.A1(G475), .A2(new_n395), .B1(new_n407), .B2(new_n410), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n521), .A2(G900), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n519), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n649), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n620), .A2(new_n525), .A3(new_n629), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT99), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n650), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n620), .A2(new_n525), .A3(new_n629), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .A4(new_n673), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n670), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XNOR2_X1  g496(.A(new_n673), .B(KEYINPUT39), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT101), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  INV_X1    g500(.A(new_n316), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n275), .B2(new_n303), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n669), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n515), .A2(new_n517), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n452), .B1(new_n396), .B2(new_n411), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n525), .A2(new_n694), .A3(new_n660), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n686), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  AOI21_X1  g512(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n408), .A2(KEYINPUT20), .A3(new_n409), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n389), .A2(KEYINPUT92), .A3(new_n354), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n390), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n702), .B2(new_n388), .ZN(new_n703));
  INV_X1    g517(.A(G475), .ZN(new_n704));
  OAI22_X1  g518(.A1(new_n699), .A2(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n617), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n679), .A2(new_n705), .A3(new_n706), .A4(new_n673), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n663), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n333), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT102), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n670), .A2(new_n712), .A3(new_n708), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  NAND2_X1  g529(.A1(new_n565), .A2(new_n568), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n559), .B1(new_n716), .B2(new_n394), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(new_n569), .ZN(new_n718));
  INV_X1    g532(.A(new_n529), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n333), .A2(new_n609), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n634), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n333), .A2(new_n609), .A3(new_n651), .A4(new_n720), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND2_X1  g540(.A1(new_n679), .A2(new_n720), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n661), .A2(new_n621), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n453), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n333), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  OAI21_X1  g545(.A(new_n317), .B1(new_n304), .B2(new_n274), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n323), .B1(new_n326), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n328), .A2(new_n317), .A3(new_n329), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n319), .B(KEYINPUT73), .ZN(new_n735));
  AOI21_X1  g549(.A(G902), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n609), .B(new_n733), .C1(new_n736), .C2(new_n637), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n720), .A2(new_n621), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n671), .A2(new_n675), .A3(KEYINPUT103), .A4(new_n452), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n695), .B2(new_n679), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  AND3_X1   g558(.A1(new_n642), .A2(new_n661), .A3(new_n733), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n708), .A2(new_n745), .A3(new_n720), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n668), .A2(new_n331), .B1(G472), .B2(new_n307), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n645), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n333), .A2(KEYINPUT105), .A3(new_n609), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n618), .A2(new_n673), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n526), .B1(new_n515), .B2(new_n517), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n570), .A2(KEYINPUT104), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n529), .C1(new_n562), .C2(new_n569), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n752), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n750), .A2(new_n751), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n673), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n671), .A2(new_n617), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n333), .A2(new_n609), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n758), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR2_X1   g581(.A1(new_n650), .A2(new_n761), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n333), .A2(new_n609), .A3(new_n768), .A4(new_n763), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NOR2_X1   g584(.A1(new_n557), .A2(new_n547), .ZN(new_n771));
  INV_X1    g585(.A(new_n548), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT45), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n773), .B2(KEYINPUT45), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n560), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  INV_X1    g592(.A(new_n569), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n529), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n683), .A3(new_n753), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n671), .A2(new_n706), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT43), .Z(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n644), .A3(new_n661), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n785), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NAND4_X1  g606(.A1(new_n749), .A2(new_n762), .A3(new_n645), .A4(new_n753), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n782), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n341), .ZN(G42));
  NOR2_X1   g612(.A1(new_n650), .A2(new_n528), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n640), .A2(new_n799), .A3(new_n643), .A4(new_n652), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n725), .B(new_n800), .C1(new_n634), .C2(new_n721), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n743), .A2(new_n730), .A3(new_n665), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n745), .A2(new_n762), .A3(new_n763), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n514), .A2(KEYINPUT86), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n511), .B1(new_n628), .B2(new_n492), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n517), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n525), .B(new_n673), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n453), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n333), .A2(new_n709), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n769), .A2(new_n804), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n765), .B2(new_n760), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n671), .A2(new_n528), .A3(new_n617), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n640), .A2(new_n814), .A3(new_n643), .A4(new_n652), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n610), .A2(new_n815), .A3(KEYINPUT106), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT106), .B1(new_n610), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n803), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n712), .B1(new_n670), .B2(new_n708), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n749), .A2(new_n707), .A3(KEYINPUT102), .A4(new_n663), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n681), .B(new_n746), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n740), .A2(new_n742), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT107), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n660), .B2(new_n673), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n606), .A2(KEYINPUT107), .A3(new_n658), .A4(new_n761), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n662), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT108), .B(new_n662), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n823), .A2(new_n831), .A3(new_n690), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n822), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n822), .B2(new_n832), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(KEYINPUT109), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n822), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n823), .A2(new_n831), .A3(new_n690), .ZN(new_n838));
  AND4_X1   g652(.A1(KEYINPUT109), .A2(new_n837), .A3(KEYINPUT52), .A4(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(KEYINPUT53), .B(new_n819), .C1(new_n836), .C2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n681), .A2(new_n746), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n714), .A3(new_n838), .A4(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n819), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g662(.A(KEYINPUT110), .B(KEYINPUT53), .C1(new_n845), .C2(new_n819), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n840), .B(new_n841), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n819), .B1(new_n836), .B2(new_n839), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n847), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n803), .A2(new_n813), .A3(new_n818), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n844), .B2(new_n835), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n841), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n787), .A2(new_n520), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n737), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n794), .A2(new_n796), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n718), .A2(new_n529), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n753), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n720), .A2(new_n753), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n690), .A2(new_n864), .A3(new_n645), .A4(new_n519), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n671), .A3(new_n617), .ZN(new_n866));
  INV_X1    g680(.A(new_n745), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n859), .A2(new_n864), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n863), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n526), .A2(new_n860), .A3(new_n693), .A4(new_n720), .ZN(new_n870));
  NOR2_X1   g684(.A1(KEYINPUT111), .A2(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n869), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n869), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n750), .A2(new_n751), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT48), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n859), .A2(new_n727), .A3(new_n737), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n865), .A2(new_n618), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(G952), .A3(new_n335), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n881), .A2(new_n883), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n858), .A2(new_n876), .A3(new_n877), .A4(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(G952), .A2(G953), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n718), .B(KEYINPUT49), .Z(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n609), .A3(new_n525), .A4(new_n529), .ZN(new_n892));
  OR4_X1    g706(.A1(new_n690), .A2(new_n892), .A3(new_n694), .A4(new_n786), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(G75));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n485), .A2(new_n486), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n491), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT55), .Z(new_n902));
  AND2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n335), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  OAI21_X1  g720(.A(KEYINPUT110), .B1(new_n855), .B2(KEYINPUT53), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n846), .A2(new_n842), .A3(new_n847), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n394), .B1(new_n909), .B2(new_n840), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n910), .A2(KEYINPUT114), .A3(new_n776), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT114), .B1(new_n910), .B2(new_n776), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n841), .B1(new_n909), .B2(new_n840), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n851), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n560), .B(KEYINPUT113), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n716), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n905), .B1(new_n913), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(new_n408), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n408), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n905), .ZN(G60));
  XOR2_X1   g737(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n615), .A2(new_n394), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n613), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n850), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT116), .B1(new_n931), .B2(new_n905), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n851), .B2(new_n914), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT116), .ZN(new_n934));
  INV_X1    g748(.A(new_n905), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n613), .B1(new_n858), .B2(new_n927), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n932), .A2(new_n936), .A3(new_n937), .ZN(G63));
  XNOR2_X1  g752(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n437), .A2(new_n394), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n896), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n607), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n896), .A2(new_n657), .A3(new_n941), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(new_n935), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT118), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n943), .B(new_n945), .C1(new_n947), .C2(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n935), .A3(new_n944), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT61), .B1(new_n944), .B2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n951), .ZN(G66));
  NAND2_X1  g766(.A1(new_n803), .A2(new_n818), .ZN(new_n953));
  NAND2_X1  g767(.A1(G224), .A2(G953), .ZN(new_n954));
  OAI22_X1  g768(.A1(new_n953), .A2(G953), .B1(new_n523), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n900), .B1(G898), .B2(new_n335), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT119), .Z(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  AOI21_X1  g772(.A(new_n335), .B1(G227), .B2(G900), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n697), .A2(new_n837), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n797), .B1(new_n789), .B2(new_n790), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n685), .A2(new_n753), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n749), .A2(new_n645), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n677), .A2(new_n618), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT121), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n967), .A2(KEYINPUT121), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n335), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n255), .A2(new_n265), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n400), .B(KEYINPUT120), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n335), .A2(G900), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT124), .ZN(new_n978));
  INV_X1    g792(.A(new_n769), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n783), .A2(new_n683), .A3(new_n823), .ZN(new_n980));
  INV_X1    g794(.A(new_n878), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n963), .A2(new_n766), .A3(new_n837), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n983), .B2(new_n335), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n975), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n976), .B1(new_n985), .B2(KEYINPUT125), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n984), .A2(new_n987), .A3(new_n975), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n959), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n959), .B(KEYINPUT123), .Z(new_n990));
  NOR2_X1   g804(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n976), .A2(KEYINPUT122), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n976), .A2(KEYINPUT122), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n994), .ZN(G72));
  XNOR2_X1  g809(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n637), .A2(new_n394), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n971), .B2(new_n953), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n269), .B(KEYINPUT127), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n274), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n983), .B2(new_n953), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1001), .A2(new_n274), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n905), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n853), .A2(new_n856), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n998), .B1(new_n276), .B2(new_n316), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(G57));
endmodule


