//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n632, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  OR2_X1    g010(.A1(KEYINPUT0), .A2(G82), .ZN(new_n436));
  NAND2_X1  g011(.A1(KEYINPUT0), .A2(G82), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR3_X1   g027(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n453));
  NAND3_X1  g028(.A1(new_n453), .A2(new_n436), .A3(new_n437), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI22_X1  g037(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n456), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n461), .B2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G101), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(new_n477), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT68), .Z(G160));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT69), .Z(new_n490));
  NAND3_X1  g065(.A1(new_n472), .A2(G2105), .A3(new_n474), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  INV_X1    g068(.A(new_n475), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n490), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n491), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n506), .B2(G2104), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(G2104), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n474), .B(new_n505), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n472), .A2(KEYINPUT70), .A3(new_n474), .A4(new_n505), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(KEYINPUT4), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(G2104), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n471), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(new_n473), .A3(G138), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n478), .A2(KEYINPUT71), .A3(new_n517), .A4(new_n505), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n503), .B1(new_n513), .B2(new_n521), .ZN(G164));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT6), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(G543), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT5), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n524), .A2(new_n526), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G88), .ZN(new_n537));
  INV_X1    g112(.A(G75), .ZN(new_n538));
  OR3_X1    g113(.A1(new_n538), .A2(new_n530), .A3(KEYINPUT73), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT73), .B1(new_n538), .B2(new_n530), .ZN(new_n540));
  INV_X1    g115(.A(G62), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(new_n533), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n523), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n529), .A2(new_n537), .A3(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  NAND2_X1  g122(.A1(new_n528), .A2(G51), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n536), .A2(G89), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT7), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  AND2_X1   g128(.A1(G63), .A2(G651), .ZN(new_n554));
  AOI211_X1 g129(.A(new_n552), .B(new_n553), .C1(new_n534), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n548), .A2(new_n549), .A3(new_n555), .ZN(G286));
  INV_X1    g131(.A(G286), .ZN(G168));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G64), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n542), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(new_n544), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n524), .A2(G90), .A3(new_n526), .A4(new_n534), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n524), .A2(G52), .A3(G543), .A4(new_n526), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G171));
  XNOR2_X1  g139(.A(KEYINPUT74), .B(G43), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n524), .A2(G543), .A3(new_n526), .A4(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G81), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n566), .B1(new_n567), .B2(new_n523), .C1(new_n568), .C2(new_n535), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G188));
  NAND4_X1  g151(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n526), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT9), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n524), .A2(G91), .A3(new_n526), .A4(new_n534), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n534), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n525), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n578), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G299));
  NAND3_X1  g163(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G301));
  NAND4_X1  g164(.A1(new_n524), .A2(G49), .A3(G543), .A4(new_n526), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n524), .A2(G87), .A3(new_n526), .A4(new_n534), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n527), .B1(new_n535), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n531), .A2(new_n533), .A3(G61), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n597), .A2(new_n598), .B1(G73), .B2(G543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n534), .A2(KEYINPUT77), .A3(G61), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n523), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n542), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n544), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT78), .ZN(new_n608));
  AOI22_X1  g183(.A1(G47), .A2(new_n528), .B1(new_n536), .B2(G85), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(KEYINPUT79), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(new_n536), .A2(G92), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n542), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G651), .ZN(new_n620));
  INV_X1    g195(.A(G54), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n527), .B2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n624), .A2(new_n625), .B1(KEYINPUT80), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(KEYINPUT80), .B2(new_n626), .ZN(G284));
  OAI21_X1  g203(.A(new_n627), .B1(KEYINPUT80), .B2(new_n626), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT81), .Z(new_n631));
  INV_X1    g206(.A(G299), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G868), .ZN(G297));
  XOR2_X1   g208(.A(G297), .B(KEYINPUT82), .Z(G280));
  XNOR2_X1  g209(.A(new_n614), .B(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n635), .A2(new_n622), .ZN(new_n636));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n478), .A2(new_n482), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n492), .A2(G123), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n494), .A2(G135), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n473), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n667), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2084), .B(G2090), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT17), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n682), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(G2096), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n690), .A3(new_n693), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n698), .C1(new_n690), .C2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(KEYINPUT20), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT86), .Z(new_n703));
  XOR2_X1   g278(.A(G1991), .B(G1996), .Z(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n701), .B(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G21), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G168), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1966), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT31), .B(G11), .Z(new_n714));
  INV_X1    g289(.A(G28), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT30), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT94), .Z(new_n717));
  AOI21_X1  g292(.A(G29), .B1(new_n715), .B2(KEYINPUT30), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n651), .B2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(G29), .A2(G33), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n494), .A2(G139), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n482), .A2(G103), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT25), .Z(new_n725));
  AOI22_X1  g300(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n725), .C1(new_n473), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n722), .B1(new_n727), .B2(new_n720), .ZN(new_n728));
  INV_X1    g303(.A(G2072), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n721), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n713), .B(new_n730), .C1(new_n729), .C2(new_n728), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G160), .B2(new_n720), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2084), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G4), .A2(G16), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT89), .Z(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n624), .B2(new_n709), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n720), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n720), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2078), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  NAND2_X1  g323(.A1(G162), .A2(G29), .ZN(new_n749));
  OR2_X1    g324(.A1(G29), .A2(G35), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G5), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G171), .B2(G16), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1961), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n709), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n570), .B2(new_n709), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G1341), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(G1341), .ZN(new_n761));
  AND4_X1   g336(.A1(new_n754), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n738), .A2(new_n747), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G32), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n767), .A2(new_n768), .B1(new_n482), .B2(G105), .ZN(new_n769));
  INV_X1    g344(.A(G129), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n491), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G141), .B2(new_n494), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT92), .Z(new_n773));
  AOI21_X1  g348(.A(new_n764), .B1(new_n773), .B2(G29), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT93), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(KEYINPUT93), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n720), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n784));
  INV_X1    g359(.A(G140), .ZN(new_n785));
  INV_X1    g360(.A(G128), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n784), .B1(new_n475), .B2(new_n785), .C1(new_n786), .C2(new_n491), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT90), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT90), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n790), .A2(KEYINPUT91), .A3(G29), .ZN(new_n791));
  AOI21_X1  g366(.A(KEYINPUT91), .B1(new_n790), .B2(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n782), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n763), .A2(new_n780), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n709), .A2(G20), .ZN(new_n796));
  NAND2_X1  g371(.A1(G299), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(KEYINPUT23), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n798), .A2(G1956), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(G1956), .B1(new_n798), .B2(new_n800), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n752), .A2(new_n753), .A3(new_n748), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n795), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n709), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n709), .ZN(new_n809));
  INV_X1    g384(.A(G1971), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G6), .A2(G16), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n602), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G23), .ZN(new_n816));
  INV_X1    g391(.A(G288), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT33), .B(G1976), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n811), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n720), .A2(G25), .ZN(new_n825));
  OR2_X1    g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n827));
  INV_X1    g402(.A(G131), .ZN(new_n828));
  INV_X1    g403(.A(G119), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n827), .B1(new_n475), .B2(new_n828), .C1(new_n829), .C2(new_n491), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n720), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n709), .A2(G24), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G290), .B2(G16), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(G1986), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(G1986), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT87), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n821), .A2(new_n822), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n824), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT88), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n844), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n842), .ZN(new_n850));
  INV_X1    g425(.A(new_n847), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n824), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n807), .B1(new_n848), .B2(new_n852), .ZN(G311));
  OR3_X1    g428(.A1(new_n763), .A2(new_n780), .A3(new_n794), .ZN(new_n854));
  INV_X1    g429(.A(new_n806), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n851), .B1(new_n850), .B2(new_n824), .ZN(new_n858));
  AOI211_X1 g433(.A(new_n823), .B(new_n847), .C1(new_n849), .C2(new_n842), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(G150));
  NAND2_X1  g435(.A1(new_n636), .A2(G559), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n524), .A2(G93), .A3(new_n526), .A4(new_n534), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n864), .B1(new_n865), .B2(new_n523), .C1(new_n866), .C2(new_n527), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n569), .B(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n868), .B2(new_n863), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(G860), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT97), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n772), .B(KEYINPUT92), .ZN(new_n875));
  MUX2_X1   g450(.A(new_n875), .B(new_n772), .S(new_n727), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n513), .A2(new_n521), .ZN(new_n877));
  INV_X1    g452(.A(new_n503), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n790), .B(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n494), .A2(G142), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n473), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(G130), .B2(new_n492), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n644), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n831), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n881), .A2(new_n890), .A3(new_n882), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT98), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT98), .ZN(new_n895));
  XNOR2_X1  g470(.A(G160), .B(new_n496), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n651), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n892), .A2(new_n893), .ZN(new_n900));
  INV_X1    g475(.A(new_n897), .ZN(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(G395));
  AND2_X1   g482(.A1(new_n584), .A2(new_n585), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n584), .A2(new_n585), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n624), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n586), .A2(new_n636), .A3(new_n587), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n639), .B(new_n868), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT99), .B1(new_n910), .B2(new_n911), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(G290), .A2(new_n817), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n611), .A2(G288), .A3(new_n612), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G166), .A2(G305), .ZN(new_n930));
  NAND2_X1  g505(.A1(G303), .A2(new_n602), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n930), .A2(KEYINPUT100), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n930), .A2(new_n931), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(KEYINPUT100), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n927), .B(new_n928), .C1(new_n936), .C2(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n919), .A2(KEYINPUT42), .A3(new_n923), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n926), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n926), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n867), .A2(new_n625), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  XNOR2_X1  g521(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n950));
  NAND2_X1  g525(.A1(G171), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G301), .A2(KEYINPUT102), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G286), .ZN(new_n954));
  NAND3_X1  g529(.A1(G168), .A2(new_n952), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n569), .B(new_n867), .Z(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n868), .A2(new_n955), .A3(new_n954), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT103), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n956), .B2(new_n957), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n948), .A2(new_n949), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n959), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n963), .B(new_n938), .C1(new_n912), .C2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n958), .A2(new_n959), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n948), .B2(KEYINPUT104), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n913), .A2(new_n970), .A3(new_n915), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n962), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(new_n961), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n973), .B(new_n974), .C1(new_n921), .C2(new_n922), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n938), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n967), .A2(new_n976), .A3(KEYINPUT43), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n912), .A2(new_n964), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n973), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n916), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n938), .ZN(new_n982));
  INV_X1    g557(.A(new_n963), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n939), .B1(new_n983), .B2(new_n979), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n947), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n967), .B2(new_n976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n978), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(KEYINPUT44), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(G397));
  AND2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NOR2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  OR3_X1    g567(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT106), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G164), .B2(G1384), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G40), .ZN(new_n998));
  NOR4_X1   g573(.A1(new_n477), .A2(new_n481), .A3(new_n998), .A4(new_n485), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G290), .A2(KEYINPUT106), .A3(G1986), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n993), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n790), .A2(G2067), .ZN(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n788), .A2(new_n1005), .A3(new_n789), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(KEYINPUT108), .A3(new_n1006), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1000), .B1(new_n1011), .B2(new_n772), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(G1996), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n830), .A2(new_n833), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n830), .A2(new_n833), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1001), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT107), .B1(new_n1000), .B2(G1996), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1000), .A2(KEYINPUT107), .A3(G1996), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n773), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AND4_X1   g596(.A1(new_n1003), .A2(new_n1014), .A3(new_n1017), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n584), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT57), .A4(new_n583), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1956), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  INV_X1    g606(.A(G1384), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n519), .A2(new_n520), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n517), .B1(new_n509), .B2(new_n510), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n512), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1031), .B(new_n1032), .C1(new_n1035), .C2(new_n503), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n999), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n879), .B2(new_n1032), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1030), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT45), .B(new_n1032), .C1(new_n1035), .C2(new_n503), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT56), .B(G2072), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n996), .A2(new_n1043), .A3(new_n999), .A4(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1029), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT120), .B(new_n1029), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1032), .B(new_n1039), .C1(new_n1035), .C2(new_n503), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1052), .A2(new_n999), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n879), .A2(new_n1032), .A3(new_n999), .ZN(new_n1055));
  OAI22_X1  g630(.A1(new_n1054), .A2(G1348), .B1(G2067), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n636), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1051), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1041), .A2(new_n1059), .A3(new_n1045), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n624), .A2(KEYINPUT122), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n624), .A2(KEYINPUT122), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(new_n1067), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT121), .B(G1996), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n996), .A2(new_n1043), .A3(new_n999), .A4(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n1055), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT59), .B1(new_n1073), .B2(new_n570), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n1075), .B(new_n569), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1059), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1060), .B1(new_n1078), .B2(KEYINPUT61), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1041), .A2(new_n1059), .A3(new_n1080), .A4(new_n1045), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1058), .A2(new_n1060), .B1(new_n1068), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT45), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(G164), .B2(G1384), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1032), .B(new_n994), .C1(new_n1035), .C2(new_n503), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n999), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  OR3_X1    g663(.A1(new_n1087), .A2(new_n1088), .A3(G2078), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1052), .A2(new_n999), .A3(new_n1053), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT125), .B(G1961), .Z(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n996), .A2(new_n1093), .A3(new_n1043), .A4(new_n999), .ZN(new_n1094));
  AOI21_X1  g669(.A(G171), .B1(new_n1094), .B2(new_n1088), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT126), .B1(new_n1094), .B2(new_n1088), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1094), .A2(new_n1088), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1092), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1094), .A2(KEYINPUT126), .A3(new_n1088), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(G301), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1094), .A2(new_n1088), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1089), .A2(new_n1104), .A3(new_n1092), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT54), .B1(new_n1105), .B2(G171), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1102), .A2(KEYINPUT54), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1087), .A2(new_n712), .ZN(new_n1108));
  INV_X1    g683(.A(G2084), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1052), .A2(new_n1109), .A3(new_n1053), .A4(new_n999), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(G168), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT124), .B1(new_n1111), .B2(G8), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT51), .B1(new_n1112), .B2(KEYINPUT123), .ZN(new_n1113));
  OR2_X1    g688(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1054), .A2(new_n1109), .B1(new_n1087), .B2(new_n712), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(G168), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G286), .A2(KEYINPUT124), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n590), .A2(new_n591), .A3(G1976), .A4(new_n592), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT111), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(new_n1055), .A3(G8), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT52), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT112), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT113), .B(G1976), .Z(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(G288), .B2(new_n1129), .ZN(new_n1130));
  AND4_X1   g705(.A1(G8), .A2(new_n1122), .A3(new_n1055), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1055), .A2(G8), .ZN(new_n1132));
  INV_X1    g707(.A(new_n596), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n1134));
  INV_X1    g709(.A(new_n601), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(G1981), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(G1981), .B1(new_n601), .B2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n601), .B2(new_n596), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1138), .A3(KEYINPUT115), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1132), .B1(KEYINPUT49), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT49), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1136), .A2(new_n1138), .A3(KEYINPUT115), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1131), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n996), .A2(new_n1043), .A3(new_n999), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n810), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1090), .A2(G2090), .ZN(new_n1147));
  OAI21_X1  g722(.A(G8), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(G303), .A2(G8), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT55), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(KEYINPUT110), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1128), .B(new_n1143), .C1(new_n1148), .C2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1145), .B1(new_n1158), .B2(G2090), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1155), .B1(new_n1159), .B2(G8), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1120), .A2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1083), .A2(new_n1107), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(G8), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1054), .A2(new_n748), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1145), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1156), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n1167), .B2(new_n1166), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1128), .A2(new_n1143), .ZN(new_n1170));
  NAND2_X1  g745(.A1(G168), .A2(G8), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1115), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT63), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  OR3_X1    g749(.A1(new_n1115), .A2(KEYINPUT63), .A3(new_n1171), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1175), .A2(new_n1160), .B1(new_n1156), .B2(new_n1148), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G305), .A2(G1981), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G288), .A2(G1976), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1132), .B1(new_n1180), .B2(KEYINPUT116), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT116), .ZN(new_n1182));
  AOI211_X1 g757(.A(G1976), .B(G288), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(new_n1177), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1176), .A2(new_n1170), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1105), .A2(G171), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1157), .A2(new_n1186), .A3(new_n1160), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1113), .A2(new_n1119), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1174), .B(new_n1185), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1022), .B1(new_n1163), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1019), .A2(KEYINPUT46), .A3(new_n1020), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT46), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1020), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(new_n1018), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1012), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT47), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1014), .A2(new_n1016), .A3(new_n1021), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1000), .B1(new_n1200), .B2(new_n1006), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n992), .A2(new_n1001), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT48), .ZN(new_n1203));
  AND4_X1   g778(.A1(new_n1017), .A2(new_n1014), .A3(new_n1021), .A4(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1199), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1193), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(new_n977), .A2(new_n985), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n466), .A2(G227), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n673), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n673), .A2(new_n1209), .A3(KEYINPUT127), .ZN(new_n1213));
  AOI21_X1  g787(.A(G229), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g788(.A(new_n902), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n894), .A2(new_n898), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n1214), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1208), .A2(new_n1217), .ZN(G308));
  OAI211_X1 g792(.A(new_n903), .B(new_n1214), .C1(new_n985), .C2(new_n977), .ZN(G225));
endmodule


