//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n206), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n217), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G226), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n253), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n262), .A2(KEYINPUT70), .A3(G226), .A4(new_n259), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n255), .A2(new_n257), .A3(G232), .A4(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n252), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT66), .A2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n270), .B(G274), .C1(new_n275), .C2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G238), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n252), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n250), .B1(new_n269), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n270), .A2(G274), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT66), .A2(G41), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT66), .A2(G41), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n279), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G238), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n267), .B1(new_n261), .B2(new_n263), .ZN(new_n290));
  OAI211_X1 g0090(.A(KEYINPUT13), .B(new_n289), .C1(new_n290), .C2(new_n252), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT14), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n281), .A2(new_n291), .A3(new_n292), .A4(G169), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n281), .A2(new_n291), .A3(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT14), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n269), .A2(new_n280), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n269), .B2(new_n280), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n203), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n256), .A2(G20), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n311));
  INV_X1    g0111(.A(G50), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n225), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(KEYINPUT11), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n270), .B2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n309), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT11), .B1(new_n315), .B2(new_n317), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n305), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n300), .A2(new_n301), .A3(G190), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n281), .A2(G200), .A3(new_n291), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT8), .B(G58), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT67), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n202), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n310), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n314), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n317), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n306), .A2(G50), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n319), .B2(G50), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(KEYINPUT9), .A3(new_n344), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G222), .A2(G1698), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n259), .A2(G223), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n262), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n352), .C1(G77), .C2(new_n262), .ZN(new_n353));
  INV_X1    g0153(.A(G226), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n276), .C1(new_n354), .C2(new_n279), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G200), .B2(new_n355), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n347), .A2(new_n348), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT10), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n345), .B(new_n362), .C1(G179), .C2(new_n355), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n276), .B1(new_n212), .B2(new_n279), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n262), .A2(G232), .A3(new_n259), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n262), .A2(G238), .A3(G1698), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n365), .B(new_n366), .C1(new_n213), .C2(new_n262), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n364), .B1(new_n352), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n317), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT68), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n310), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n332), .A2(new_n314), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G20), .B2(G77), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n371), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n319), .A2(G77), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G77), .B2(new_n306), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n370), .B1(G169), .B2(new_n368), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n377), .A2(new_n379), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n368), .A2(G190), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n368), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT69), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n331), .A2(new_n360), .A3(new_n363), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n262), .B2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n203), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n204), .A2(new_n205), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n313), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n388), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT73), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n254), .A3(G33), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n401), .A3(new_n257), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n402), .A2(new_n389), .A3(new_n226), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n389), .B1(new_n402), .B2(new_n226), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(new_n203), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n313), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n398), .B(new_n317), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n354), .B2(G1698), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(new_n399), .A3(new_n257), .A4(new_n401), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n252), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n252), .A2(G232), .A3(new_n278), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n276), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n383), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n354), .A2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G223), .B2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n412), .B1(new_n402), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n352), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n252), .A2(G232), .A3(new_n278), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT74), .B1(new_n287), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n276), .A2(new_n423), .A3(new_n414), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n420), .A2(new_n422), .A3(new_n424), .A4(new_n356), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n336), .A2(new_n319), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n336), .B2(new_n306), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n408), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT76), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT76), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n408), .A2(new_n426), .A3(new_n432), .A4(new_n429), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n408), .A2(new_n426), .A3(new_n435), .A4(new_n429), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT77), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n431), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n433), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n398), .A2(new_n317), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n404), .A2(new_n203), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n402), .A2(new_n389), .A3(new_n226), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n407), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n429), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n361), .B1(new_n413), .B2(new_n415), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n420), .A2(new_n422), .A3(new_n424), .A4(new_n369), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n446), .B1(new_n445), .B2(new_n450), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT75), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT7), .B1(new_n258), .B2(new_n226), .ZN(new_n455));
  AOI211_X1 g0255(.A(new_n389), .B(G20), .C1(new_n255), .C2(new_n257), .ZN(new_n456));
  OAI21_X1  g0256(.A(G68), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n406), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n371), .B1(new_n458), .B2(new_n388), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n399), .A2(new_n401), .A3(new_n257), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT7), .B1(new_n460), .B2(G20), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G68), .A3(new_n443), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n428), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT18), .B1(new_n464), .B2(new_n449), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n454), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n439), .B(new_n440), .C1(new_n453), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n387), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n214), .A2(G1698), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G257), .B2(G1698), .ZN(new_n472));
  INV_X1    g0272(.A(G303), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n402), .A2(new_n472), .B1(new_n473), .B2(new_n262), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n352), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n270), .B(G45), .C1(new_n476), .C2(G41), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n283), .B2(new_n284), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(G274), .A4(new_n252), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT5), .B1(new_n273), .B2(new_n274), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n252), .B1(new_n481), .B2(new_n477), .ZN(new_n482));
  INV_X1    g0282(.A(G270), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n475), .B(new_n480), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n307), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n270), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n371), .A2(new_n306), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n316), .A2(new_n225), .B1(G20), .B2(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(new_n226), .C1(G33), .C2(new_n218), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT20), .B1(new_n489), .B2(new_n491), .ZN(new_n493));
  OAI221_X1 g0293(.A(new_n486), .B1(new_n488), .B2(new_n485), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n484), .A2(G169), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n474), .A2(new_n352), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n497), .A2(new_n498), .A3(new_n369), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n496), .B1(new_n499), .B2(new_n494), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n484), .A2(KEYINPUT21), .A3(G169), .A4(new_n494), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n498), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n361), .B1(new_n504), .B2(new_n475), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT82), .A3(KEYINPUT21), .A4(new_n494), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(G190), .A3(new_n475), .ZN(new_n507));
  INV_X1    g0307(.A(new_n494), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n497), .A2(new_n498), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n383), .C2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n500), .A2(new_n503), .A3(new_n506), .A4(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n511), .A2(KEYINPUT83), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(KEYINPUT83), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g0314(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n515));
  NOR2_X1   g0315(.A1(new_n306), .A2(G107), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n213), .B2(new_n488), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT22), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n226), .A2(G87), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n258), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n519), .A2(new_n522), .A3(G20), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(new_n399), .A3(new_n257), .A4(new_n401), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT84), .B1(new_n226), .B2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT23), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI211_X1 g0327(.A(KEYINPUT84), .B(new_n527), .C1(new_n226), .C2(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n310), .A2(G116), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n521), .A2(new_n524), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT24), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n526), .A2(new_n528), .B1(G116), .B2(new_n310), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n524), .A4(new_n521), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n518), .B1(new_n536), .B2(new_n317), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n219), .A2(G1698), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(G250), .B2(G1698), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n460), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n252), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G264), .B(new_n252), .C1(new_n481), .C2(new_n477), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n480), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G190), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n537), .B(new_n547), .C1(new_n383), .C2(new_n546), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n543), .A2(new_n545), .A3(G179), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n352), .B1(new_n478), .B2(new_n479), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n477), .B1(new_n275), .B2(new_n476), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n252), .A2(G274), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n550), .A2(G264), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n542), .B1(new_n402), .B2(new_n539), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n352), .ZN(new_n556));
  AOI21_X1  g0356(.A(G169), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n371), .B1(new_n532), .B2(new_n535), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n518), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n554), .A2(new_n369), .A3(new_n556), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n546), .B2(G169), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT86), .B1(new_n537), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n548), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G274), .ZN(new_n566));
  INV_X1    g0366(.A(G250), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(KEYINPUT79), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n286), .A2(G1), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT79), .B(G250), .C1(new_n286), .C2(G1), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n352), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n212), .A2(G1698), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G238), .B2(G1698), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n573), .B1(new_n402), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n369), .B(new_n572), .C1(new_n352), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n352), .ZN(new_n578));
  INV_X1    g0378(.A(new_n572), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n361), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT80), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G238), .A2(G1698), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n212), .B2(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n583), .A2(new_n399), .A3(new_n257), .A4(new_n401), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n252), .B1(new_n584), .B2(new_n573), .ZN(new_n585));
  OAI21_X1  g0385(.A(G169), .B1(new_n585), .B2(new_n572), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n578), .A2(G179), .A3(new_n579), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT81), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT68), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n372), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n372), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n590), .B1(new_n594), .B2(new_n488), .ZN(new_n595));
  INV_X1    g0395(.A(new_n488), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n373), .A2(new_n596), .A3(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n306), .B1(new_n592), .B2(new_n593), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n226), .B1(new_n266), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n522), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n226), .A2(G33), .A3(G97), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n601), .A2(new_n603), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n203), .A2(G20), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n399), .A2(new_n401), .A3(new_n257), .A4(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n371), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n598), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n581), .A2(new_n589), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n212), .A2(G1698), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n399), .A2(new_n401), .A3(new_n257), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT4), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n490), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G250), .A2(G1698), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n259), .A2(G244), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n614), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n262), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n352), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n219), .B(new_n352), .C1(new_n478), .C2(new_n479), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n480), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n361), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT6), .ZN(new_n627));
  AND2_X1   g0427(.A1(G97), .A2(G107), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n602), .ZN(new_n629));
  NAND2_X1  g0429(.A1(KEYINPUT6), .A2(G97), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT78), .B1(new_n630), .B2(G107), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT78), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n213), .A3(KEYINPUT6), .A4(G97), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n313), .A2(G77), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n213), .B1(new_n390), .B2(new_n391), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n317), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n306), .A2(G97), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n488), .B2(new_n218), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n621), .A2(new_n352), .B1(G257), .B2(new_n550), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(new_n369), .A3(new_n480), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n626), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(G107), .B1(new_n455), .B2(new_n456), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n634), .A2(G20), .B1(G77), .B2(new_n313), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n642), .B1(new_n650), .B2(new_n317), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n622), .A2(new_n624), .A3(G190), .A4(new_n480), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n252), .B1(new_n615), .B2(new_n620), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n552), .A2(new_n481), .A3(new_n477), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(new_n623), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n651), .B(new_n652), .C1(new_n383), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n578), .A2(new_n579), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G200), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n488), .A2(new_n522), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n599), .A2(new_n608), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n578), .A2(G190), .A3(new_n579), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n611), .A2(new_n647), .A3(new_n656), .A4(new_n662), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n470), .A2(new_n514), .A3(new_n565), .A4(new_n663), .ZN(G372));
  NAND2_X1  g0464(.A1(new_n439), .A2(new_n440), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n330), .A2(new_n380), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n326), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n451), .A2(new_n452), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n360), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n363), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n647), .A2(new_n656), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n658), .A2(new_n661), .A3(new_n660), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n577), .B2(new_n580), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n586), .A2(KEYINPUT87), .A3(new_n588), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n679), .B2(new_n610), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n674), .A2(new_n680), .A3(new_n548), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n500), .A2(new_n506), .A3(new_n503), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n537), .A2(new_n563), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(G169), .B1(new_n645), .B2(new_n480), .ZN(new_n686));
  NOR4_X1   g0486(.A1(new_n653), .A2(new_n623), .A3(G179), .A4(new_n654), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n651), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n611), .A3(new_n662), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT26), .ZN(new_n690));
  INV_X1    g0490(.A(new_n678), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT87), .B1(new_n586), .B2(new_n588), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n610), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT26), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n688), .A3(new_n694), .A4(new_n662), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n690), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT88), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n690), .A2(new_n698), .A3(new_n695), .A4(new_n693), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n685), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n673), .B1(new_n470), .B2(new_n700), .ZN(G369));
  NAND3_X1  g0501(.A1(new_n270), .A2(new_n226), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G343), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n494), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT90), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n682), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n514), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n565), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n708), .B1(new_n560), .B2(new_n518), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n683), .B2(new_n708), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n682), .A2(new_n707), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n683), .A2(new_n707), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT91), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n717), .A2(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n229), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n275), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n603), .A2(G116), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n726), .A2(new_n270), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n224), .B2(new_n726), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g0531(.A1(new_n697), .A2(new_n699), .ZN(new_n732));
  INV_X1    g0532(.A(new_n685), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n708), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n561), .A2(new_n564), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n682), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n681), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n688), .A2(new_n611), .A3(new_n694), .A4(new_n662), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n677), .A2(new_n678), .B1(new_n609), .B2(new_n598), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n647), .A3(new_n675), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n693), .B(new_n740), .C1(new_n742), .C2(new_n694), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n707), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n565), .A2(new_n663), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n707), .C1(new_n512), .C2(new_n513), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  INV_X1    g0549(.A(new_n657), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n546), .A3(new_n645), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n509), .A2(G179), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n546), .A2(G179), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(new_n484), .A3(new_n625), .A4(new_n657), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n657), .A2(new_n543), .A3(new_n545), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n499), .A4(new_n645), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n753), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n758), .B2(new_n708), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT93), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n759), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n748), .B(new_n761), .C1(new_n763), .C2(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G330), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n746), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n731), .B1(new_n766), .B2(G1), .ZN(G364));
  AOI21_X1  g0567(.A(new_n225), .B1(G20), .B2(new_n361), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n226), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n369), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n356), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n772), .A2(G311), .B1(G326), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n769), .B1(new_n777), .B2(G20), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n779), .A2(KEYINPUT98), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(KEYINPUT98), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n775), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT99), .Z(new_n785));
  NOR2_X1   g0585(.A1(new_n383), .A2(G179), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n769), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n262), .B1(new_n788), .B2(G283), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n773), .A2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(KEYINPUT33), .A2(G317), .ZN(new_n791));
  AND2_X1   g0591(.A1(KEYINPUT33), .A2(G317), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n226), .A2(new_n356), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n770), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n789), .B(new_n793), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n777), .A2(new_n226), .A3(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G329), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n795), .A2(new_n786), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n799), .B1(new_n803), .B2(new_n473), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n785), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n782), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G97), .ZN(new_n807));
  INV_X1    g0607(.A(new_n774), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n312), .ZN(new_n809));
  INV_X1    g0609(.A(new_n790), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n262), .B1(new_n787), .B2(new_n213), .C1(new_n810), .C2(new_n203), .ZN(new_n811));
  INV_X1    g0611(.A(new_n803), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n809), .B(new_n811), .C1(new_n812), .C2(G87), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n798), .A2(G159), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT32), .Z(new_n815));
  OAI22_X1  g0615(.A1(new_n796), .A2(new_n202), .B1(new_n771), .B2(new_n211), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT95), .ZN(new_n817));
  AND4_X1   g0617(.A1(new_n807), .A2(new_n813), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n768), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n226), .A2(G13), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n270), .B1(new_n820), .B2(G45), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n726), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n724), .A2(new_n258), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(G355), .B1(new_n485), .B2(new_n724), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n248), .A2(new_n286), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n460), .A2(new_n724), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(G45), .B2(new_n223), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(G13), .A2(G33), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(G20), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n768), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT94), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n824), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n833), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n819), .B(new_n837), .C1(new_n712), .C2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT100), .Z(new_n840));
  NOR2_X1   g0640(.A1(new_n712), .A2(G330), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n713), .A2(new_n824), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(G396));
  INV_X1    g0643(.A(new_n768), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n832), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n823), .B1(G77), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n810), .A2(new_n847), .B1(new_n808), .B2(new_n473), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n796), .A2(new_n783), .B1(new_n771), .B2(new_n485), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n258), .B1(new_n787), .B2(new_n522), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n812), .A2(G107), .B1(G311), .B2(new_n798), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n807), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n460), .B1(new_n203), .B2(new_n787), .C1(new_n803), .C2(new_n312), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G132), .B2(new_n798), .ZN(new_n855));
  INV_X1    g0655(.A(new_n796), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n856), .A2(G143), .B1(new_n772), .B2(G159), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n774), .A2(G137), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n340), .C2(new_n810), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n855), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n782), .A2(new_n202), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n846), .B1(new_n865), .B2(new_n768), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n384), .B1(new_n381), .B2(new_n707), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n380), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n380), .A2(new_n708), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n870), .B2(new_n832), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n734), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n700), .A2(new_n385), .A3(new_n708), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n765), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n824), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n872), .A2(new_n765), .A3(new_n873), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT101), .Z(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G384));
  OR2_X1    g0679(.A1(new_n634), .A2(KEYINPUT35), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n634), .A2(KEYINPUT35), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(G116), .A3(new_n227), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT36), .Z(new_n883));
  NAND3_X1  g0683(.A1(new_n224), .A2(G77), .A3(new_n393), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n312), .A2(G68), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n270), .B(G13), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n324), .B(new_n708), .C1(new_n305), .C2(new_n330), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n324), .A2(new_n708), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n303), .B1(new_n294), .B2(new_n295), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n329), .B(new_n889), .C1(new_n890), .C2(new_n323), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n869), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n317), .B1(new_n405), .B2(new_n407), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n462), .B2(new_n406), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n429), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n706), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n468), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n706), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n464), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT37), .B1(new_n445), .B2(new_n450), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(new_n431), .A3(new_n433), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n449), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n431), .A2(new_n906), .A3(new_n433), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT102), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT37), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(new_n907), .B2(KEYINPUT37), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n899), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT103), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n468), .B2(new_n898), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(KEYINPUT103), .A3(new_n911), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n912), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n894), .A2(new_n919), .B1(new_n669), .B2(new_n706), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n922), .B1(new_n669), .B2(new_n706), .C1(new_n894), .C2(new_n919), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n439), .A2(new_n669), .A3(new_n440), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n901), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n430), .B1(new_n464), .B2(new_n449), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n926), .B2(new_n901), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n904), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n913), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n919), .B2(new_n932), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n326), .A2(new_n707), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n921), .A2(new_n923), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n746), .A2(new_n470), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n672), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n938), .B(new_n940), .Z(new_n941));
  INV_X1    g0741(.A(G330), .ZN(new_n942));
  INV_X1    g0742(.A(new_n912), .ZN(new_n943));
  AND4_X1   g0743(.A1(KEYINPUT103), .A2(new_n899), .A3(KEYINPUT38), .A4(new_n911), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT103), .B1(new_n917), .B2(new_n911), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n748), .A2(new_n763), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n947), .A2(new_n870), .A3(new_n892), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n931), .A2(new_n913), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n948), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n946), .A2(new_n950), .B1(new_n952), .B2(KEYINPUT40), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n469), .A2(new_n947), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n942), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n941), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n270), .B2(new_n820), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n941), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n887), .B1(new_n959), .B2(new_n960), .ZN(G367));
  OR3_X1    g0761(.A1(new_n693), .A2(new_n660), .A3(new_n707), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n680), .B1(new_n660), .B2(new_n707), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n674), .B1(new_n651), .B2(new_n707), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n688), .A2(new_n708), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n719), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT42), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n969), .B(KEYINPUT107), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n561), .A2(new_n564), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n647), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n972), .B1(new_n707), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n966), .B(new_n976), .C1(KEYINPUT43), .C2(new_n964), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n966), .ZN(new_n978));
  INV_X1    g0778(.A(new_n717), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(new_n973), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n978), .B(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n726), .B(KEYINPUT41), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n722), .A2(new_n970), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT44), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n722), .A2(new_n970), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n716), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n719), .B1(new_n989), .B2(new_n718), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n713), .B(new_n990), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n766), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n979), .B1(new_n984), .B2(new_n986), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n982), .B1(new_n994), .B2(new_n766), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n981), .B1(new_n995), .B2(new_n822), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n806), .A2(G68), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n772), .A2(G50), .B1(G159), .B2(new_n790), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT110), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n262), .B1(new_n787), .B2(new_n211), .C1(new_n340), .C2(new_n796), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G143), .B2(new_n774), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n812), .A2(G58), .B1(G137), .B2(new_n798), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n782), .A2(new_n213), .B1(new_n847), .B2(new_n771), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT109), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n812), .A2(G116), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT46), .ZN(new_n1007));
  INV_X1    g0807(.A(G311), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n810), .A2(new_n783), .B1(new_n808), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n788), .A2(G97), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1010), .B(new_n402), .C1(new_n473), .C2(new_n796), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G317), .C2(new_n798), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1003), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT47), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n844), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n237), .A2(new_n828), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n835), .B1(new_n724), .B2(new_n373), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n824), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT108), .Z(new_n1021));
  OAI211_X1 g0821(.A(new_n1017), .B(new_n1021), .C1(new_n838), .C2(new_n964), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n996), .A2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n991), .A2(new_n822), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n728), .A2(new_n825), .B1(new_n213), .B2(new_n724), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n241), .A2(new_n286), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n332), .A2(G50), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT50), .Z(new_n1028));
  OAI211_X1 g0828(.A(new_n727), .B(new_n286), .C1(new_n203), .C2(new_n211), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n828), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1025), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n824), .B1(new_n1031), .B2(new_n836), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n782), .A2(new_n594), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G150), .A2(new_n798), .B1(new_n337), .B2(new_n790), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n211), .B2(new_n803), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1010), .B1(new_n312), .B2(new_n796), .C1(new_n203), .C2(new_n771), .ZN(new_n1036));
  INV_X1    g0836(.A(G159), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n460), .B1(new_n808), .B2(new_n1037), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n856), .A2(G317), .B1(new_n772), .B2(G303), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n808), .B2(new_n794), .C1(new_n1008), .C2(new_n810), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1041), .A2(new_n1042), .B1(new_n783), .B2(new_n803), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G283), .B2(new_n806), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n798), .A2(G326), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n402), .C1(new_n485), .C2(new_n787), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1046), .B2(KEYINPUT49), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1039), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1032), .B1(new_n989), .B2(new_n838), .C1(new_n1051), .C2(new_n844), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n992), .A2(new_n726), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n766), .A2(new_n991), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1024), .B(new_n1052), .C1(new_n1053), .C2(new_n1054), .ZN(G393));
  OAI21_X1  g0855(.A(new_n992), .B1(new_n988), .B2(new_n993), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n994), .A2(new_n726), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT115), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n994), .A2(KEYINPUT115), .A3(new_n726), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n988), .A2(new_n821), .A3(new_n993), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n973), .A2(new_n833), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n772), .A2(G294), .B1(G303), .B2(new_n790), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n782), .B2(new_n485), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT113), .Z(new_n1066));
  AOI22_X1  g0866(.A1(new_n856), .A2(G311), .B1(G317), .B2(new_n774), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n798), .A2(G322), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n258), .B1(new_n213), .B2(new_n787), .C1(new_n803), .C2(new_n847), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n812), .A2(G68), .B1(G143), .B2(new_n798), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n808), .A2(new_n340), .B1(new_n796), .B2(new_n1037), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n332), .A2(new_n771), .B1(new_n787), .B2(new_n522), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n402), .B(new_n1075), .C1(G50), .C2(new_n790), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G77), .B2(new_n806), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n768), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n828), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n836), .B1(new_n218), .B2(new_n229), .C1(new_n245), .C2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT112), .Z(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n823), .A3(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT114), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1062), .B1(new_n1063), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1061), .A2(new_n1085), .ZN(G390));
  AOI21_X1  g0886(.A(new_n942), .B1(new_n748), .B2(new_n763), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n469), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n673), .B(new_n1088), .C1(new_n746), .C2(new_n470), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n385), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n734), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n869), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n765), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n892), .B1(new_n1094), .B2(new_n870), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n892), .A2(new_n870), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1087), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1093), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1094), .A2(new_n870), .A3(new_n892), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n707), .B(new_n868), .C1(new_n739), .C2(new_n743), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT116), .B1(new_n1101), .B2(new_n869), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n869), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1087), .A2(new_n870), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1100), .B(new_n1105), .C1(new_n892), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1099), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1090), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n946), .A2(KEYINPUT39), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n893), .B1(new_n734), .B2(new_n1091), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n892), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n935), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1113), .A3(new_n933), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n935), .B(new_n951), .C1(new_n1105), .C2(new_n1112), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(new_n1100), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1097), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(KEYINPUT117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n869), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1119), .A2(new_n1102), .A3(new_n1112), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n951), .A2(new_n935), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n931), .A2(new_n932), .A3(new_n913), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n946), .B2(KEYINPUT39), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n1124), .B2(new_n1113), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1097), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1109), .B1(new_n1118), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1125), .B2(new_n1097), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n936), .B1(new_n1093), .B2(new_n892), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1115), .B1(new_n934), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(KEYINPUT117), .A3(new_n1098), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1089), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1129), .A2(new_n1132), .A3(new_n1116), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n726), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1129), .A2(new_n1132), .A3(new_n822), .A4(new_n1116), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n823), .B1(new_n337), .B2(new_n845), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n803), .A2(new_n340), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n856), .A2(G132), .B1(new_n772), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n258), .B1(new_n788), .B2(G50), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n790), .A2(G137), .B1(new_n774), .B2(G128), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G125), .B2(new_n798), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1139), .B(new_n1146), .C1(new_n1037), .C2(new_n782), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n812), .A2(G87), .B1(G294), .B2(new_n798), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n810), .A2(new_n213), .B1(new_n808), .B2(new_n847), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n796), .A2(new_n485), .B1(new_n771), .B2(new_n218), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n258), .B1(new_n787), .B2(new_n203), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1149), .B(new_n1153), .C1(new_n782), .C2(new_n211), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1148), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1137), .B1(new_n1156), .B2(new_n768), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n934), .B2(new_n832), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT119), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1136), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1135), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT120), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT120), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1135), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(G378));
  NAND2_X1  g0965(.A1(new_n1134), .A2(new_n1090), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n360), .A2(new_n363), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n900), .B1(new_n342), .B2(new_n344), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OR3_X1    g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n953), .B2(new_n942), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n948), .A2(new_n949), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n919), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n949), .B1(new_n951), .B2(new_n948), .ZN(new_n1181));
  OAI211_X1 g0981(.A(G330), .B(new_n1176), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n938), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n920), .A2(KEYINPUT104), .B1(new_n934), .B2(new_n936), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1185), .A2(new_n1178), .A3(new_n923), .A4(new_n1182), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1167), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1166), .A2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1134), .A2(new_n1090), .B1(new_n1186), .B2(new_n1184), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1188), .B(new_n726), .C1(KEYINPUT57), .C2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n823), .B1(G50), .B2(new_n845), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n312), .B1(G33), .B2(G41), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n402), .B2(new_n285), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n856), .A2(G107), .B1(new_n788), .B2(G58), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n485), .B2(new_n808), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G97), .B2(new_n790), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n460), .B(new_n275), .C1(new_n812), .C2(G77), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n798), .A2(G283), .B1(new_n373), .B2(new_n772), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n997), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT58), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n803), .A2(new_n1140), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n856), .A2(G128), .B1(new_n772), .B2(G137), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n774), .A2(G125), .ZN(new_n1204));
  INV_X1    g1004(.A(G132), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1204), .C1(new_n1205), .C2(new_n810), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1202), .B(new_n1206), .C1(new_n806), .C2(G150), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n256), .B(new_n272), .C1(new_n787), .C2(new_n1037), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n798), .B2(G124), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT59), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1201), .B1(new_n1200), .B2(new_n1199), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1191), .B1(new_n1214), .B2(new_n768), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1176), .B2(new_n832), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n822), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1190), .A2(new_n1219), .ZN(G375));
  NOR2_X1   g1020(.A1(new_n1133), .A2(new_n982), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1090), .B2(new_n1108), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT121), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1112), .A2(new_n831), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n823), .B1(G68), .B2(new_n845), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n202), .A2(new_n787), .B1(new_n771), .B2(new_n340), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n402), .B(new_n1226), .C1(new_n798), .C2(G128), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n1037), .B2(new_n803), .C1(new_n782), .C2(new_n312), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT122), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n856), .A2(G137), .B1(new_n1141), .B2(new_n790), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1205), .B2(new_n808), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n810), .A2(new_n485), .B1(new_n808), .B2(new_n783), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n796), .A2(new_n847), .B1(new_n771), .B2(new_n213), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n258), .B1(new_n787), .B2(new_n211), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n798), .A2(G303), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n218), .C2(new_n803), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1229), .A2(new_n1231), .B1(new_n1033), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1225), .B1(new_n1238), .B2(new_n768), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1108), .A2(new_n822), .B1(new_n1224), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1223), .A2(new_n1240), .ZN(G381));
  OR4_X1    g1041(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n996), .A2(new_n1061), .A3(new_n1022), .A4(new_n1085), .ZN(new_n1243));
  OR4_X1    g1043(.A1(new_n1161), .A2(new_n1242), .A3(G375), .A4(new_n1243), .ZN(G407));
  INV_X1    g1044(.A(G375), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1161), .ZN(new_n1246));
  INV_X1    g1046(.A(G343), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G213), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(G407), .A2(G213), .A3(new_n1250), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1090), .B2(new_n1108), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1089), .A2(KEYINPUT60), .A3(new_n1099), .A4(new_n1107), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1255), .A2(new_n726), .A3(new_n1109), .A4(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n878), .A3(new_n1240), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n878), .B1(new_n1257), .B2(new_n1240), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1240), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(G384), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(KEYINPUT124), .A3(new_n1258), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1249), .A2(G2897), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1261), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT125), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT125), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1261), .A2(new_n1264), .A3(new_n1268), .A4(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1263), .A2(new_n1258), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1270), .A2(new_n1265), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1162), .A2(new_n1164), .A3(new_n1190), .A4(new_n1219), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1218), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1184), .A2(KEYINPUT123), .A3(new_n1186), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n822), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1189), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1277), .B(new_n1216), .C1(new_n1278), .C2(new_n982), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1246), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1249), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1252), .B1(new_n1272), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1243), .ZN(new_n1285));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1285), .B(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1273), .A2(new_n1280), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n1248), .A3(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1291), .A2(KEYINPUT63), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(KEYINPUT63), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1283), .B(new_n1288), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1261), .A2(KEYINPUT62), .A3(new_n1264), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1281), .A2(new_n1296), .ZN(new_n1297));
  XOR2_X1   g1097(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1298));
  AOI22_X1  g1098(.A1(new_n1295), .A2(new_n1297), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1281), .A2(KEYINPUT127), .A3(new_n1296), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1282), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1294), .B1(new_n1301), .B2(new_n1288), .ZN(G405));
  INV_X1    g1102(.A(new_n1273), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1246), .B2(G375), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1270), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1290), .B2(new_n1304), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1288), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1285), .B(new_n1286), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1308), .B(new_n1305), .C1(new_n1290), .C2(new_n1304), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(G402));
endmodule


