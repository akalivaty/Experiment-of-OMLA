//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G134), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT11), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n197), .A3(G134), .ZN(new_n202));
  AOI211_X1 g016(.A(G131), .B(new_n198), .C1(new_n200), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n202), .ZN(new_n205));
  INV_X1    g019(.A(new_n198), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n196), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT2), .A2(G113), .ZN(new_n209));
  NAND3_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G116), .B(G119), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT2), .A2(G113), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n209), .A3(new_n214), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n188), .A2(new_n190), .A3(new_n224), .A4(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n187), .A2(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n225), .B(new_n227), .C1(G128), .C2(new_n193), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n201), .B1(G134), .B2(new_n197), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n199), .A2(KEYINPUT11), .A3(G137), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n204), .B(new_n206), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n197), .B2(G134), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n199), .A3(G137), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n197), .A2(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n228), .A2(new_n231), .A3(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n208), .A2(new_n223), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G237), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G237), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT68), .B(G953), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G210), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT27), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n244), .A2(new_n245), .A3(new_n248), .A4(G210), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n239), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n237), .A2(new_n231), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n237), .A2(new_n231), .A3(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n228), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT30), .B1(new_n261), .B2(new_n208), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n208), .A2(KEYINPUT30), .A3(new_n238), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n222), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n256), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g080(.A(new_n207), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n195), .B1(new_n267), .B2(new_n231), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n188), .A2(new_n190), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n269), .A2(new_n270), .B1(KEYINPUT1), .B2(new_n226), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n257), .A2(new_n258), .B1(new_n271), .B2(new_n225), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n272), .B2(new_n260), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n222), .B(new_n263), .C1(new_n273), .C2(KEYINPUT30), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n256), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n266), .A2(KEYINPUT31), .A3(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n273), .A2(new_n223), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n239), .A2(KEYINPUT28), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n239), .A2(KEYINPUT28), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n255), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT70), .B1(new_n265), .B2(KEYINPUT31), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n274), .A2(new_n284), .A3(new_n285), .A4(new_n256), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n277), .A2(new_n282), .A3(new_n283), .A4(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n283), .A2(new_n286), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(KEYINPUT71), .A3(new_n282), .A4(new_n277), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT72), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n239), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n274), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n255), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n255), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n278), .A2(new_n280), .A3(new_n303), .A4(new_n279), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n223), .B1(new_n208), .B2(new_n238), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n239), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n310), .A2(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n255), .A2(new_n305), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT73), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n294), .B1(new_n289), .B2(new_n291), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n298), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G217), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(G234), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n245), .A2(G221), .A3(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G137), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n270), .A2(G119), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n270), .A2(KEYINPUT23), .A3(G119), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n330), .A2(G128), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n335), .B(new_n331), .C1(new_n336), .C2(KEYINPUT23), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n338));
  INV_X1    g152(.A(G110), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n337), .B2(KEYINPUT75), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n334), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G125), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT16), .ZN(new_n346));
  OR3_X1    g160(.A1(new_n344), .A2(KEYINPUT16), .A3(G140), .ZN(new_n347));
  AOI21_X1  g161(.A(G146), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n347), .A3(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n350), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n348), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n332), .A2(new_n333), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n337), .B2(G110), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n343), .A2(new_n345), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n187), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n351), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n328), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n360), .A3(new_n328), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n323), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n355), .A2(new_n360), .A3(new_n328), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(new_n361), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n325), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n324), .A2(G902), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n370), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n376), .A2(new_n379), .A3(new_n383), .A4(new_n380), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n386), .A3(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n222), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n375), .A2(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n378), .A2(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(G101), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n214), .A2(KEYINPUT5), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n330), .A3(G116), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n395), .A2(new_n330), .A3(KEYINPUT80), .A4(G116), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(G113), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n393), .A2(new_n400), .A3(new_n221), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n388), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n388), .A2(new_n403), .A3(new_n401), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n195), .A2(G125), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(KEYINPUT81), .C1(G125), .C2(new_n228), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n271), .A2(new_n410), .A3(new_n344), .A4(new_n225), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G953), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G224), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT82), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n402), .A2(new_n420), .A3(new_n404), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n407), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(KEYINPUT7), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n409), .A2(new_n411), .A3(new_n423), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n406), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n403), .B(KEYINPUT8), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n400), .A2(new_n221), .B1(new_n384), .B2(new_n391), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(KEYINPUT83), .B2(new_n401), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n393), .A2(new_n400), .A3(new_n432), .A4(new_n221), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n323), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n374), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n407), .A2(new_n419), .A3(new_n421), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n439));
  INV_X1    g253(.A(new_n430), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n433), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n428), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(new_n406), .A3(new_n426), .A4(new_n425), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n438), .A2(new_n443), .A3(new_n323), .A4(new_n373), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n437), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n443), .A3(new_n323), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT84), .A3(new_n374), .ZN(new_n447));
  NAND2_X1  g261(.A1(G234), .A2(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G952), .A3(new_n413), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT90), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n245), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(G902), .A3(new_n448), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT91), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n445), .A2(new_n447), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n352), .A2(new_n354), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n244), .A2(new_n245), .A3(G214), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT85), .B(G143), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n189), .A2(KEYINPUT85), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n244), .A2(new_n245), .A3(G214), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G131), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n204), .A3(new_n468), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n204), .B1(new_n466), .B2(new_n468), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT17), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n474), .B2(KEYINPUT17), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n463), .B(new_n473), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G113), .B(G122), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(new_n375), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n358), .A2(new_n187), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n359), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n469), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n469), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n469), .B2(new_n484), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n478), .A2(new_n480), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n480), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n469), .A2(new_n484), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n485), .B1(new_n495), .B2(new_n488), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n466), .A2(new_n204), .A3(new_n468), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n474), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n358), .B(KEYINPUT19), .Z(new_n499));
  OAI21_X1  g313(.A(new_n351), .B1(new_n499), .B2(G146), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n493), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G475), .A2(G902), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n462), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  AOI211_X1 g320(.A(KEYINPUT20), .B(new_n506), .C1(new_n492), .C2(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n478), .A2(new_n491), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n493), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n509), .B2(new_n492), .ZN(new_n510));
  INV_X1    g324(.A(G475), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n505), .A2(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT13), .B1(new_n270), .B2(G143), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n199), .ZN(new_n514));
  XNOR2_X1  g328(.A(G128), .B(G143), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G116), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT88), .ZN(new_n519));
  INV_X1    g333(.A(G116), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G122), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(new_n378), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n378), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n518), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n521), .B(KEYINPUT14), .ZN(new_n527));
  OAI21_X1  g341(.A(G107), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n519), .A2(new_n378), .A3(new_n521), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n515), .B(new_n199), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT9), .B(G234), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n533), .A2(new_n322), .A3(G953), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n531), .A3(new_n534), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G478), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n540), .B(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n512), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G221), .B1(new_n533), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G469), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n245), .A2(G227), .ZN(new_n548));
  XOR2_X1   g362(.A(G110), .B(G140), .Z(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n225), .A2(KEYINPUT77), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT77), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n193), .A2(new_n553), .A3(new_n224), .A4(G128), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n271), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n393), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n203), .A2(new_n207), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n385), .A2(new_n196), .A3(new_n387), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n393), .A2(KEYINPUT10), .A3(new_n228), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n558), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n556), .B1(new_n228), .B2(new_n393), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT78), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n564), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n559), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n563), .B2(new_n567), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n551), .B(new_n562), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n567), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n551), .B1(new_n572), .B2(new_n562), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n570), .B1(new_n573), .B2(KEYINPUT79), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT79), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n575), .B(new_n551), .C1(new_n572), .C2(new_n562), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n547), .B(new_n323), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n547), .A2(new_n323), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n562), .B1(new_n568), .B2(new_n569), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n562), .A2(new_n551), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n579), .A2(new_n550), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n581), .B2(G469), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n546), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n461), .A2(new_n544), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n461), .A2(new_n544), .A3(KEYINPUT92), .A4(new_n583), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n321), .A2(new_n372), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT93), .B(G101), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G3));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT33), .B1(new_n534), .B2(KEYINPUT95), .ZN(new_n592));
  INV_X1    g406(.A(new_n537), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n534), .B1(new_n524), .B2(new_n531), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n592), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n536), .A2(new_n537), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n541), .A2(G902), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n591), .A2(new_n595), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n595), .A2(new_n597), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n598), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(new_n538), .B2(G478), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n512), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n446), .B2(new_n374), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n458), .B1(new_n609), .B2(new_n444), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n446), .A2(KEYINPUT94), .A3(new_n374), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n456), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n292), .B2(new_n323), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n583), .A2(new_n372), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n617), .A2(new_n319), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n492), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n480), .B1(new_n478), .B2(new_n491), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n323), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G475), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n626), .B(new_n543), .C1(new_n505), .C2(new_n507), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n613), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n619), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT98), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n617), .A2(new_n319), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT25), .B1(new_n368), .B2(new_n323), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n367), .A2(new_n361), .A3(new_n365), .A4(G902), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n324), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n355), .A2(new_n360), .ZN(new_n639));
  INV_X1    g453(.A(new_n328), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n371), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n635), .A2(new_n586), .A3(new_n587), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  NAND2_X1  g461(.A1(new_n609), .A2(new_n444), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(new_n644), .A3(new_n611), .A4(new_n457), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n577), .A2(new_n582), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n545), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n451), .B1(new_n453), .B2(new_n652), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n649), .A2(new_n651), .A3(new_n627), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n318), .B1(new_n319), .B2(KEYINPUT32), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n297), .B(new_n294), .C1(new_n289), .C2(new_n291), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT99), .B(G128), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G30));
  NAND2_X1  g473(.A1(new_n445), .A2(new_n447), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT100), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n660), .B(new_n662), .Z(new_n663));
  XOR2_X1   g477(.A(new_n653), .B(KEYINPUT39), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n583), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n512), .A2(new_n543), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n458), .A3(new_n644), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n616), .B1(new_n310), .B2(new_n255), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n266), .A2(new_n276), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(G472), .A2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT102), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n319), .B2(KEYINPUT32), .ZN(new_n675));
  OAI221_X1 g489(.A(new_n669), .B1(KEYINPUT40), .B2(new_n665), .C1(new_n656), .C2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT103), .B(G143), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G45));
  INV_X1    g492(.A(new_n653), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n512), .A2(new_n604), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n649), .A2(new_n680), .A3(new_n651), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n655), .B2(new_n656), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(G146), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G48));
  NOR2_X1   g498(.A1(new_n547), .A2(KEYINPUT105), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n574), .A2(new_n576), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n685), .B1(new_n686), .B2(G902), .ZN(new_n687));
  OAI221_X1 g501(.A(new_n323), .B1(KEYINPUT105), .B2(new_n547), .C1(new_n574), .C2(new_n576), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n545), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n372), .B(new_n690), .C1(new_n655), .C2(new_n656), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n614), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT41), .B(G113), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NOR2_X1   g508(.A1(new_n691), .A2(new_n629), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n520), .ZN(G18));
  NOR3_X1   g510(.A1(new_n512), .A2(new_n456), .A3(new_n543), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n689), .A2(new_n649), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n697), .B(new_n698), .C1(new_n655), .C2(new_n656), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  NAND2_X1  g514(.A1(new_n292), .A2(new_n323), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT106), .A3(G472), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  AOI21_X1  g517(.A(G902), .B1(new_n289), .B2(new_n291), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n703), .B1(new_n704), .B2(new_n616), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n290), .B(new_n277), .C1(new_n303), .C2(new_n313), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n702), .A2(new_n705), .B1(new_n295), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n610), .A2(new_n512), .A3(new_n543), .A4(new_n611), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n456), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n372), .A3(new_n690), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n295), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n649), .A2(new_n689), .A3(new_n680), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT106), .B1(new_n701), .B2(G472), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n704), .A2(new_n703), .A3(new_n616), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n712), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  NAND2_X1  g531(.A1(new_n320), .A2(KEYINPUT108), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n656), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n718), .A2(new_n720), .A3(new_n298), .A4(new_n318), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT107), .B1(new_n660), .B2(new_n457), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n723), .B(new_n458), .C1(new_n445), .C2(new_n447), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n722), .A2(new_n724), .A3(new_n680), .A4(new_n651), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n721), .A2(KEYINPUT42), .A3(new_n372), .A4(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n722), .A2(new_n724), .A3(new_n651), .ZN(new_n728));
  INV_X1    g542(.A(new_n680), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n372), .B1(new_n655), .B2(new_n656), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  INV_X1    g548(.A(new_n372), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n627), .A3(new_n653), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n321), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  INV_X1    g552(.A(new_n722), .ZN(new_n739));
  INV_X1    g553(.A(new_n724), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n579), .A2(new_n550), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n580), .A2(new_n572), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n547), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n581), .A2(KEYINPUT45), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n578), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n577), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(KEYINPUT109), .A3(new_n545), .A4(new_n664), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n545), .B1(new_n749), .B2(new_n750), .ZN(new_n754));
  INV_X1    g568(.A(new_n664), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n741), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n512), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n604), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n601), .A2(new_n603), .ZN(new_n761));
  INV_X1    g575(.A(new_n599), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n763), .B2(new_n512), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n296), .B1(new_n616), .B2(new_n704), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n644), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT44), .A4(new_n644), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n757), .B(new_n769), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  NOR4_X1   g589(.A1(new_n321), .A2(new_n372), .A3(new_n680), .A4(new_n741), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n545), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n754), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NAND3_X1  g596(.A1(new_n760), .A2(new_n451), .A3(new_n764), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT115), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n372), .A3(new_n690), .A4(new_n707), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n612), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n721), .A2(new_n372), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n741), .A2(new_n689), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT117), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n787), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n786), .B1(new_n793), .B2(KEYINPUT48), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n675), .A2(new_n656), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n372), .A2(new_n788), .A3(new_n451), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n607), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n413), .A2(G952), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT118), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n787), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n784), .A2(new_n791), .A3(new_n788), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n791), .B1(new_n784), .B2(new_n788), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT48), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n783), .B(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n372), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(new_n689), .ZN(new_n810));
  INV_X1    g624(.A(new_n663), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n458), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n458), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n785), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n707), .A2(new_n644), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n802), .B2(new_n803), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n796), .A2(new_n758), .A3(new_n763), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n808), .A2(new_n809), .A3(new_n741), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n687), .A2(new_n688), .A3(new_n546), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n777), .A2(new_n779), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n819), .A2(KEYINPUT51), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n794), .B(new_n806), .C1(new_n817), .C2(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n827));
  XNOR2_X1  g641(.A(new_n822), .B(KEYINPUT116), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n821), .B1(new_n780), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n819), .A2(new_n829), .A3(new_n820), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n827), .B1(new_n830), .B2(new_n816), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n512), .A2(new_n604), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n461), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n628), .A2(new_n461), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT111), .B1(new_n605), .B2(new_n460), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT112), .B1(new_n627), .B2(new_n460), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n835), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n619), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n841), .A2(new_n645), .A3(new_n699), .ZN(new_n842));
  INV_X1    g656(.A(new_n691), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n615), .B2(new_n630), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n588), .A3(new_n844), .A4(new_n710), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n702), .A2(new_n705), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n725), .A3(new_n644), .A4(new_n712), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n638), .A2(new_n643), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n848), .A2(new_n512), .A3(new_n543), .A4(new_n653), .ZN(new_n849));
  OAI221_X1 g663(.A(new_n728), .B1(new_n736), .B2(new_n849), .C1(new_n655), .C2(new_n656), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n733), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n583), .A2(new_n848), .A3(new_n679), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n708), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n675), .B2(new_n656), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n716), .A2(new_n657), .A3(new_n682), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n707), .A2(new_n713), .B1(new_n321), .B2(new_n654), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n682), .A2(new_n857), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n862), .A4(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n858), .A2(new_n859), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n853), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n588), .A2(new_n645), .A3(new_n699), .A4(new_n841), .ZN(new_n867));
  INV_X1    g681(.A(new_n709), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n809), .A2(new_n689), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n691), .B1(new_n614), .B2(new_n629), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n847), .A2(new_n850), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n732), .B2(new_n726), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n862), .A2(KEYINPUT52), .A3(new_n657), .A4(new_n716), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  AND4_X1   g689(.A1(KEYINPUT53), .A2(new_n871), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT54), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n875), .A3(new_n873), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n871), .A4(new_n873), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n832), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n735), .A2(new_n458), .A3(new_n546), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n758), .A3(new_n604), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n687), .A2(new_n688), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n795), .A3(new_n811), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n885), .A2(new_n892), .ZN(G75));
  NAND2_X1  g707(.A1(new_n880), .A2(new_n881), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(G210), .A3(G902), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n407), .A2(new_n421), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n419), .ZN(new_n898));
  XOR2_X1   g712(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n245), .A2(G952), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G51));
  XNOR2_X1  g718(.A(new_n578), .B(KEYINPUT57), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n880), .A2(new_n882), .A3(new_n881), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n882), .B1(new_n880), .B2(new_n881), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n686), .B(KEYINPUT120), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n894), .A2(G902), .A3(new_n747), .A4(new_n746), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n903), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND2_X1  g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT121), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n894), .A2(G902), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n503), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n903), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n600), .B(new_n921), .C1(new_n906), .C2(new_n907), .ZN(new_n922));
  INV_X1    g736(.A(new_n903), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n600), .B1(new_n884), .B2(new_n921), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n880), .B2(new_n881), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(new_n368), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n642), .B(KEYINPUT122), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n930), .A2(KEYINPUT61), .A3(new_n923), .A4(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n923), .B1(new_n929), .B2(new_n368), .ZN(new_n935));
  INV_X1    g749(.A(new_n928), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n894), .A2(new_n936), .A3(new_n931), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n934), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n933), .A2(new_n938), .ZN(G66));
  INV_X1    g753(.A(G224), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n455), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n871), .B2(new_n452), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n897), .B1(G898), .B2(new_n245), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  AOI21_X1  g759(.A(new_n245), .B1(G227), .B2(G900), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT125), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n263), .B1(new_n273), .B2(KEYINPUT30), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n499), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n676), .A2(new_n682), .A3(new_n861), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n833), .A2(new_n628), .ZN(new_n955));
  OR4_X1    g769(.A1(new_n731), .A2(new_n665), .A3(new_n741), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n774), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n954), .B1(new_n774), .B2(new_n956), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n953), .B(new_n781), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n960), .B2(new_n245), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n452), .A2(G900), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n781), .A2(new_n737), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n708), .B1(new_n752), .B2(new_n756), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n801), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n733), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n774), .A2(new_n682), .A3(new_n861), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n963), .B1(new_n969), .B2(new_n245), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n948), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n774), .A2(new_n956), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n974));
  AOI22_X1  g788(.A1(new_n974), .A2(new_n957), .B1(new_n780), .B2(new_n776), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n452), .B1(new_n975), .B2(new_n953), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n972), .B(new_n947), .C1(new_n976), .C2(new_n950), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n977), .ZN(G72));
  XOR2_X1   g792(.A(new_n672), .B(KEYINPUT63), .Z(new_n979));
  NOR2_X1   g793(.A1(new_n302), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n266), .B(new_n276), .C1(new_n301), .C2(new_n981), .ZN(new_n982));
  OAI221_X1 g796(.A(new_n979), .B1(new_n980), .B2(new_n982), .C1(new_n866), .C2(new_n876), .ZN(new_n983));
  INV_X1    g797(.A(new_n979), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n969), .B2(new_n871), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n274), .A2(new_n255), .A3(new_n299), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT126), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n983), .B(new_n923), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n300), .A2(new_n303), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n975), .A2(new_n871), .A3(new_n953), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n979), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n988), .A2(new_n991), .ZN(G57));
endmodule


