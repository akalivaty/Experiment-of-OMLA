//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G15gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G22gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G15gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT88), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(G15gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n202), .A2(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n206), .A2(new_n211), .B1(KEYINPUT16), .B2(new_n207), .ZN(new_n214));
  OAI21_X1  g013(.A(G8gat), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT89), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT90), .B(G8gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n212), .B(new_n218), .C1(new_n214), .C2(KEYINPUT89), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT14), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT15), .A4(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n228), .A2(new_n229), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n231), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n238));
  INV_X1    g037(.A(new_n236), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n230), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n237), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT91), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n215), .B(new_n240), .C1(new_n217), .C2(new_n219), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT92), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n254));
  INV_X1    g053(.A(new_n211), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n210), .B1(new_n208), .B2(new_n209), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(new_n216), .A3(new_n212), .A4(new_n218), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n215), .A4(new_n240), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(new_n262), .A3(new_n245), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n247), .B(KEYINPUT13), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n248), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G141gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G197gat), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT11), .B(G169gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n270), .B(KEYINPUT12), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n251), .A2(new_n265), .A3(new_n266), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n265), .A2(KEYINPUT93), .A3(new_n266), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n251), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT93), .B1(new_n265), .B2(new_n266), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT94), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT94), .B(new_n271), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G127gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G127gat), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n291), .A2(new_n293), .A3(G134gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n290), .B2(G134gat), .ZN(new_n296));
  INV_X1    g095(.A(G134gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n289), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n287), .A2(new_n301), .A3(new_n288), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT25), .B1(new_n305), .B2(G169gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND3_X1  g119(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(G190gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT67), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n325), .A3(KEYINPUT67), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT64), .B(G169gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n305), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n320), .ZN(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n333), .B(new_n334), .C1(G183gat), .C2(G190gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n327), .A2(new_n328), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT27), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(G190gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT28), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT27), .B(G183gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n309), .A2(new_n349), .A3(new_n310), .ZN(new_n350));
  NOR2_X1   g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n351), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT68), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT68), .B1(new_n350), .B2(new_n352), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n303), .B1(new_n337), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G227gat), .ZN(new_n357));
  INV_X1    g156(.A(G233gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n360));
  AND3_X1   g159(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT24), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n334), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n311), .A2(KEYINPUT23), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n310), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n306), .B1(new_n309), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n328), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n336), .A2(new_n329), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n300), .A2(new_n302), .ZN(new_n373));
  INV_X1    g172(.A(new_n354), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT68), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n344), .A4(new_n347), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n356), .A2(new_n359), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n356), .A2(KEYINPUT71), .A3(new_n359), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT32), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n373), .B1(new_n372), .B2(new_n376), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n384), .A2(new_n385), .B1(new_n357), .B2(new_n358), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT34), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT34), .ZN(new_n388));
  OAI221_X1 g187(.A(new_n388), .B1(new_n357), .B2(new_n358), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT33), .B1(new_n380), .B2(new_n381), .ZN(new_n391));
  XOR2_X1   g190(.A(G15gat), .B(G43gat), .Z(new_n392));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n390), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n389), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n384), .A2(new_n385), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT71), .B1(new_n399), .B2(new_n359), .ZN(new_n400));
  INV_X1    g199(.A(new_n381), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n383), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G228gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(new_n358), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(G197gat), .B(G204gat), .ZN(new_n412));
  INV_X1    g211(.A(G218gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  INV_X1    g213(.A(G211gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n411), .B(new_n412), .C1(new_n418), .C2(KEYINPUT22), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n422));
  OAI21_X1  g221(.A(G218gat), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT22), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n411), .B1(new_n425), .B2(new_n412), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G141gat), .B(G148gat), .Z(new_n429));
  INV_X1    g228(.A(G155gat), .ZN(new_n430));
  INV_X1    g229(.A(G162gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT2), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G141gat), .B(G148gat), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n433), .B(new_n432), .C1(new_n437), .C2(KEYINPUT2), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n428), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n438), .ZN(new_n444));
  INV_X1    g243(.A(new_n411), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n416), .A2(new_n417), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT22), .B1(new_n446), .B2(G218gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n412), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT29), .B1(new_n449), .B2(new_n419), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n439), .B1(new_n450), .B2(KEYINPUT81), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n441), .B1(new_n420), .B2(new_n426), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n444), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n436), .A2(new_n438), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT3), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT82), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n410), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n427), .A2(KEYINPUT80), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n441), .B1(new_n449), .B2(KEYINPUT80), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n439), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n444), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI211_X1 g269(.A(new_n409), .B(new_n443), .C1(new_n466), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT31), .B(G50gat), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n463), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  INV_X1    g273(.A(new_n443), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n461), .B2(KEYINPUT82), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n455), .A2(new_n456), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n409), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n466), .A2(new_n470), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n410), .A3(new_n475), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n407), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n390), .B1(new_n391), .B2(new_n395), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n402), .A2(new_n397), .A3(new_n394), .ZN(new_n484));
  INV_X1    g283(.A(new_n383), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n472), .B1(new_n463), .B2(new_n471), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(new_n480), .A3(new_n474), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n406), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n404), .A2(new_n482), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G1gat), .B(G29gat), .Z(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G57gat), .B(G85gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n373), .A2(new_n444), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n300), .A2(new_n438), .A3(new_n436), .A4(new_n302), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n303), .A2(new_n468), .A3(new_n469), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n497), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n458), .A2(new_n506), .A3(new_n300), .A4(new_n302), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT77), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n444), .A2(KEYINPUT3), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n440), .A3(new_n373), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n499), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n502), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n511), .A2(new_n515), .A3(new_n499), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n303), .A2(new_n468), .A3(new_n506), .A4(new_n469), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n495), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n509), .A2(new_n513), .ZN(new_n523));
  INV_X1    g322(.A(new_n502), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n495), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(new_n517), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n528), .A3(new_n515), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n503), .A2(KEYINPUT4), .B1(new_n507), .B2(KEYINPUT77), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n512), .B1(new_n530), .B2(new_n505), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n531), .B2(new_n502), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT79), .A3(new_n495), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n522), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(KEYINPUT6), .A3(new_n495), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G8gat), .B(G36gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G64gat), .B(G92gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n372), .A2(new_n376), .ZN(new_n540));
  NAND2_X1  g339(.A1(G226gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n541), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT29), .B1(new_n372), .B2(new_n376), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n543), .B(new_n428), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n441), .ZN(new_n547));
  INV_X1    g346(.A(new_n542), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n547), .A2(new_n548), .B1(new_n540), .B2(new_n544), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n539), .B(new_n546), .C1(new_n549), .C2(new_n428), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT75), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n546), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n355), .B1(new_n371), .B2(new_n370), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n548), .B1(new_n557), .B2(KEYINPUT29), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n544), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n428), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT74), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n542), .B2(new_n545), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n427), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n546), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n539), .ZN(new_n567));
  INV_X1    g366(.A(new_n550), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n566), .A2(new_n567), .B1(new_n568), .B2(KEYINPUT30), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n536), .A2(new_n555), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT35), .B1(new_n490), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT87), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(KEYINPUT87), .B(KEYINPUT35), .C1(new_n490), .C2(new_n570), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT6), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n526), .B(new_n529), .C1(new_n531), .C2(new_n502), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n520), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT35), .B1(new_n577), .B2(new_n535), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n555), .A3(new_n569), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT86), .B1(new_n490), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n578), .A2(new_n555), .A3(new_n569), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n485), .B1(new_n483), .B2(new_n484), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n487), .A2(new_n406), .A3(new_n488), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n406), .B1(new_n487), .B2(new_n488), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT86), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n581), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n580), .A4(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n563), .A2(new_n564), .A3(new_n546), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n564), .B1(new_n563), .B2(new_n546), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n567), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n568), .A2(KEYINPUT30), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n550), .A2(KEYINPUT75), .A3(new_n551), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n593), .B(new_n594), .C1(new_n552), .C2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n499), .B1(new_n528), .B2(new_n511), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT39), .B1(new_n498), .B2(new_n500), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n495), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(KEYINPUT40), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT84), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n601), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT40), .B1(new_n605), .B2(KEYINPUT83), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(KEYINPUT83), .B2(new_n605), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n596), .A2(new_n520), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n563), .A2(new_n546), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n567), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n562), .B2(new_n428), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n543), .B(new_n427), .C1(new_n544), .C2(new_n545), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT38), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n568), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n561), .B2(new_n565), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT38), .B1(new_n619), .B2(new_n612), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n618), .A2(new_n620), .A3(new_n535), .A4(new_n577), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n608), .A2(new_n621), .A3(new_n587), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n582), .B2(new_n583), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n404), .A2(KEYINPUT36), .A3(new_n486), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n535), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT79), .B1(new_n532), .B2(new_n495), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n576), .A2(new_n575), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n630), .B2(new_n533), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n596), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n622), .B(new_n626), .C1(new_n587), .C2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n282), .B1(new_n590), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT9), .ZN(new_n635));
  INV_X1    g434(.A(G71gat), .ZN(new_n636));
  INV_X1    g435(.A(G78gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT95), .ZN(new_n639));
  XOR2_X1   g438(.A(G57gat), .B(G64gat), .Z(new_n640));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n641), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G71gat), .B(G78gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n639), .A2(new_n640), .A3(new_n644), .A4(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G127gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n650), .B(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n290), .ZN(new_n655));
  XOR2_X1   g454(.A(G183gat), .B(G211gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n653), .B2(new_n655), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n648), .A2(new_n649), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n220), .A2(KEYINPUT96), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT96), .B1(new_n220), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n430), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n664), .A2(new_n666), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n659), .A2(new_n660), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n660), .ZN(new_n671));
  INV_X1    g470(.A(new_n669), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n658), .A4(new_n667), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(G99gat), .B(G106gat), .Z(new_n675));
  NAND2_X1  g474(.A1(G85gat), .A2(G92gat), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT7), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G99gat), .A2(G106gat), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n679), .A2(KEYINPUT8), .ZN(new_n680));
  NOR2_X1   g479(.A1(G85gat), .A2(G92gat), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT97), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(G85gat), .ZN(new_n683));
  INV_X1    g482(.A(G92gat), .ZN(new_n684));
  AOI22_X1  g483(.A1(KEYINPUT8), .A2(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n675), .B(new_n678), .C1(new_n682), .C2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n675), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n682), .A2(new_n687), .ZN(new_n690));
  INV_X1    g489(.A(new_n678), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n243), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n237), .ZN(new_n695));
  NAND3_X1  g494(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(G190gat), .B(G218gat), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(G134gat), .B(G162gat), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n698), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n693), .A2(new_n703), .A3(new_n695), .A4(new_n696), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n699), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n699), .B2(new_n704), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n674), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(G230gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n358), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n646), .A2(new_n647), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n690), .A2(new_n689), .A3(new_n691), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n681), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n685), .A2(new_n686), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n691), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n675), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n689), .A2(KEYINPUT98), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n712), .A2(new_n713), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT10), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n646), .A3(new_n647), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n692), .B2(new_n688), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n694), .A2(KEYINPUT10), .A3(new_n712), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n711), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n711), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n719), .B2(new_n722), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(G120gat), .B(G148gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(G176gat), .B(G204gat), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n731), .B(new_n732), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n729), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n726), .A2(new_n730), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n733), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n725), .B2(new_n728), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n709), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n634), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n536), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n207), .ZN(G1324gat));
  NAND3_X1  g541(.A1(new_n634), .A2(new_n596), .A3(new_n739), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(G8gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT16), .B(G8gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT42), .B2(new_n746), .ZN(G1325gat));
  NOR3_X1   g547(.A1(new_n740), .A2(new_n202), .A3(new_n626), .ZN(new_n749));
  INV_X1    g548(.A(new_n584), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n202), .B1(new_n740), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT100), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(G1326gat));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n587), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT43), .B(G22gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1327gat));
  NAND3_X1  g557(.A1(new_n574), .A2(new_n580), .A3(new_n589), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n632), .A2(new_n584), .A3(new_n587), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT87), .B1(new_n760), .B2(KEYINPUT35), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n633), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n707), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n674), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(KEYINPUT101), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(KEYINPUT101), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n771), .A2(new_n282), .A3(new_n738), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n767), .A2(new_n631), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT102), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n222), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  INV_X1    g575(.A(new_n707), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n768), .A2(new_n738), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n634), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n222), .A3(new_n631), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n776), .A2(new_n782), .ZN(G1328gat));
  INV_X1    g582(.A(new_n596), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(G36gat), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n779), .A2(KEYINPUT103), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT103), .B1(new_n779), .B2(new_n786), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n767), .A2(new_n596), .A3(new_n772), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(G36gat), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1329gat));
  INV_X1    g595(.A(new_n626), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n765), .A2(new_n797), .A3(new_n766), .A4(new_n772), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n750), .A2(G43gat), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n798), .A2(G43gat), .B1(new_n780), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(KEYINPUT105), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1330gat));
  INV_X1    g602(.A(new_n587), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n767), .A2(new_n804), .A3(new_n772), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G50gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n780), .A2(KEYINPUT106), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT106), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n779), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n587), .A2(G50gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT48), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n806), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n806), .B2(new_n811), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1331gat));
  NAND2_X1  g614(.A1(new_n282), .A2(new_n708), .ZN(new_n816));
  INV_X1    g615(.A(new_n738), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT107), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(new_n762), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n631), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g621(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT108), .ZN(new_n825));
  NOR2_X1   g624(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n825), .B(new_n826), .ZN(G1333gat));
  AOI21_X1  g626(.A(new_n636), .B1(new_n820), .B2(new_n797), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n750), .A2(G71gat), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n830), .B(new_n831), .ZN(G1334gat));
  NAND2_X1  g631(.A1(new_n820), .A2(new_n804), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g633(.A1(new_n282), .A2(new_n674), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT110), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n738), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n767), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n631), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n762), .A2(new_n707), .A3(new_n836), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n707), .A4(new_n836), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(KEYINPUT111), .A3(new_n841), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n631), .A2(new_n683), .A3(new_n738), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n839), .A2(new_n683), .B1(new_n847), .B2(new_n848), .ZN(G1336gat));
  NAND4_X1  g648(.A1(new_n765), .A2(new_n596), .A3(new_n766), .A4(new_n837), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(new_n850), .B2(G92gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n784), .A2(G92gat), .A3(new_n817), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n845), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(G92gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n842), .A2(new_n844), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n852), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT112), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n851), .A2(new_n853), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n862));
  AOI22_X1  g661(.A1(G92gat), .A2(new_n850), .B1(new_n857), .B2(new_n852), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n861), .B(new_n862), .C1(new_n855), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1337gat));
  INV_X1    g664(.A(G99gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n767), .A2(new_n797), .A3(new_n837), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n584), .A2(new_n866), .A3(new_n738), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n847), .B2(new_n871), .ZN(G1338gat));
  NAND4_X1  g671(.A1(new_n765), .A2(new_n804), .A3(new_n766), .A4(new_n837), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G106gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT114), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n587), .A2(G106gat), .A3(new_n817), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT115), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n879), .A3(G106gat), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n875), .A2(new_n878), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n884));
  XNOR2_X1  g683(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n885));
  INV_X1    g684(.A(new_n876), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n874), .B(new_n885), .C1(new_n847), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(G1339gat));
  NOR2_X1   g687(.A1(new_n263), .A2(new_n264), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n248), .B1(new_n244), .B2(new_n245), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n270), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n738), .A2(new_n273), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n723), .A2(new_n711), .A3(new_n724), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n894), .A2(new_n725), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n711), .B(new_n898), .C1(new_n723), .C2(new_n724), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT119), .B1(new_n899), .B2(new_n733), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n723), .A2(new_n724), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n727), .A3(new_n897), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(new_n736), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n896), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n893), .B1(new_n905), .B2(KEYINPUT55), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n894), .A2(new_n725), .A3(new_n895), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n733), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n903), .B1(new_n902), .B2(new_n736), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT55), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(KEYINPUT120), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n735), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n905), .B2(KEYINPUT55), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n892), .B1(new_n916), .B2(new_n282), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n777), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n707), .A2(new_n273), .A3(new_n891), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n913), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n771), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n282), .A2(new_n708), .A3(new_n817), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT117), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n282), .A2(new_n708), .A3(new_n927), .A4(new_n817), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n536), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n490), .A2(new_n596), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n282), .ZN(new_n933));
  AOI21_X1  g732(.A(G113gat), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n804), .B1(new_n924), .B2(new_n929), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n631), .A3(new_n784), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n750), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n282), .A2(new_n285), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(G1340gat));
  AOI21_X1  g738(.A(G120gat), .B1(new_n932), .B2(new_n738), .ZN(new_n940));
  INV_X1    g739(.A(new_n936), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n750), .A2(new_n283), .A3(new_n817), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1341gat));
  NAND2_X1  g742(.A1(new_n291), .A2(new_n293), .ZN(new_n944));
  INV_X1    g743(.A(new_n937), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n923), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n932), .A2(new_n291), .A3(new_n293), .A4(new_n768), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1342gat));
  AND3_X1   g747(.A1(new_n932), .A2(new_n297), .A3(new_n707), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G134gat), .B1(new_n945), .B2(new_n777), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G1343gat));
  NOR2_X1   g753(.A1(new_n797), .A2(new_n587), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n596), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n282), .A2(G141gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n930), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n924), .A2(new_n929), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT57), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(new_n963), .A3(new_n804), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n797), .A2(new_n536), .A3(new_n596), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n915), .B1(KEYINPUT55), .B2(new_n905), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n892), .B1(new_n282), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n920), .B1(new_n967), .B2(new_n777), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(new_n768), .ZN(new_n969));
  INV_X1    g768(.A(new_n929), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n804), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT57), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n964), .A2(new_n933), .A3(new_n965), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n961), .B1(new_n973), .B2(G141gat), .ZN(new_n974));
  NOR2_X1   g773(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n974), .B(new_n975), .ZN(G1344gat));
  AND2_X1   g775(.A1(new_n930), .A2(new_n957), .ZN(new_n977));
  INV_X1    g776(.A(G148gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n978), .A3(new_n738), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT122), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n972), .ZN(new_n981));
  AOI211_X1 g780(.A(KEYINPUT59), .B(new_n978), .C1(new_n981), .C2(new_n738), .ZN(new_n982));
  XNOR2_X1  g781(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n771), .B1(new_n918), .B2(new_n921), .ZN(new_n984));
  OAI211_X1 g783(.A(KEYINPUT57), .B(new_n804), .C1(new_n984), .C2(new_n970), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n925), .B1(new_n968), .B2(new_n768), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT57), .B1(new_n986), .B2(new_n804), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n985), .B1(new_n987), .B2(KEYINPUT124), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n989));
  AOI211_X1 g788(.A(new_n989), .B(KEYINPUT57), .C1(new_n986), .C2(new_n804), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n738), .B(new_n965), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n983), .B1(new_n991), .B2(G148gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n980), .B1(new_n982), .B2(new_n992), .ZN(G1345gat));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n430), .A3(new_n768), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n981), .A2(new_n771), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n994), .B1(new_n995), .B2(new_n430), .ZN(G1346gat));
  AOI21_X1  g795(.A(G162gat), .B1(new_n977), .B2(new_n707), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n777), .A2(new_n431), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n981), .B2(new_n998), .ZN(G1347gat));
  NOR2_X1   g798(.A1(new_n490), .A2(new_n784), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n962), .A2(new_n536), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1001), .A2(new_n330), .A3(new_n933), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n596), .A2(new_n536), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n750), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n935), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g805(.A(G169gat), .B1(new_n1006), .B2(new_n282), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1003), .A2(new_n1007), .ZN(G1348gat));
  AOI21_X1  g807(.A(G176gat), .B1(new_n1001), .B2(new_n738), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1006), .A2(new_n304), .A3(new_n817), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1349gat));
  OAI21_X1  g810(.A(KEYINPUT126), .B1(new_n1006), .B2(new_n923), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n935), .A2(new_n1013), .A3(new_n771), .A4(new_n1005), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1012), .A2(G183gat), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1001), .A2(new_n345), .A3(new_n768), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(KEYINPUT60), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT60), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1015), .A2(new_n1019), .A3(new_n1016), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n1020), .ZN(G1350gat));
  NAND3_X1  g820(.A1(new_n1001), .A2(new_n342), .A3(new_n707), .ZN(new_n1022));
  OAI21_X1  g821(.A(G190gat), .B1(new_n1006), .B2(new_n777), .ZN(new_n1023));
  AND2_X1   g822(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1024));
  NOR2_X1   g823(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G1351gat));
  NOR2_X1   g825(.A1(new_n956), .A2(new_n784), .ZN(new_n1027));
  AND3_X1   g826(.A1(new_n962), .A2(new_n536), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n933), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n988), .A2(new_n990), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1030), .A2(new_n797), .A3(new_n1004), .ZN(new_n1031));
  AND2_X1   g830(.A1(new_n933), .A2(G197gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G1352gat));
  NOR2_X1   g832(.A1(new_n797), .A2(new_n1004), .ZN(new_n1034));
  OAI211_X1 g833(.A(new_n738), .B(new_n1034), .C1(new_n988), .C2(new_n990), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1035), .A2(G204gat), .ZN(new_n1036));
  NOR2_X1   g835(.A1(new_n817), .A2(G204gat), .ZN(new_n1037));
  NAND4_X1  g836(.A1(new_n962), .A2(new_n536), .A3(new_n1027), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g837(.A(KEYINPUT62), .ZN(new_n1039));
  XNOR2_X1  g838(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1041), .A2(KEYINPUT127), .ZN(new_n1042));
  INV_X1    g841(.A(KEYINPUT127), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1036), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n1042), .A2(new_n1044), .ZN(G1353gat));
  NAND4_X1  g844(.A1(new_n1028), .A2(new_n416), .A3(new_n417), .A4(new_n768), .ZN(new_n1046));
  OAI211_X1 g845(.A(new_n768), .B(new_n1034), .C1(new_n988), .C2(new_n990), .ZN(new_n1047));
  AND3_X1   g846(.A1(new_n1047), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1048));
  AOI21_X1  g847(.A(KEYINPUT63), .B1(new_n1047), .B2(G211gat), .ZN(new_n1049));
  OAI21_X1  g848(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(G1354gat));
  NAND3_X1  g849(.A1(new_n1028), .A2(new_n413), .A3(new_n707), .ZN(new_n1051));
  OAI211_X1 g850(.A(new_n707), .B(new_n1034), .C1(new_n988), .C2(new_n990), .ZN(new_n1052));
  INV_X1    g851(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g852(.A(new_n1051), .B1(new_n1053), .B2(new_n413), .ZN(G1355gat));
endmodule


