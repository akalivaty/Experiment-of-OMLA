//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT77), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT76), .B1(new_n192), .B2(G125), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G140), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n196), .A2(new_n199), .B1(G125), .B2(new_n192), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n195), .B1(new_n200), .B2(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n201), .B(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT75), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n211), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n203), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n212), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n205), .B2(new_n210), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n201), .A2(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n198), .A2(G140), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n193), .A3(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n220), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n191), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n218), .A2(new_n225), .ZN(new_n227));
  INV_X1    g041(.A(new_n190), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G217), .ZN(new_n230));
  INV_X1    g044(.A(G902), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(G234), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT74), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n231), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(KEYINPUT78), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT78), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n240), .B2(KEYINPUT79), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n239), .A2(new_n240), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n243), .B2(new_n233), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT0), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(new_n208), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT64), .A2(G146), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT64), .A2(G146), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n202), .A2(G143), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n208), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n202), .A2(G143), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n222), .B2(G143), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n259), .B2(new_n248), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT64), .A2(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT64), .A2(G146), .ZN(new_n262));
  OAI21_X1  g076(.A(G143), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n258), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(new_n257), .A3(new_n264), .A4(new_n248), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n256), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(G137), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n270), .A2(new_n272), .A3(new_n277), .A4(new_n273), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(KEYINPUT66), .A3(G131), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n246), .B1(new_n267), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n263), .A2(new_n283), .A3(G128), .A4(new_n264), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n252), .A2(new_n253), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n208), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n273), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n269), .A2(G137), .ZN(new_n289));
  OAI21_X1  g103(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n278), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n263), .A2(new_n264), .A3(new_n248), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n293), .A2(new_n265), .B1(new_n255), .B2(new_n254), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(KEYINPUT67), .A3(new_n280), .A4(new_n279), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n299));
  INV_X1    g113(.A(G113), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT68), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT2), .A3(G113), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n301), .A2(new_n303), .B1(new_n299), .B2(new_n300), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(G116), .B2(new_n206), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT69), .B(G116), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n206), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G116), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n306), .A3(G119), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n309), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n206), .A2(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n314), .B2(G119), .ZN(new_n319));
  AOI211_X1 g133(.A(KEYINPUT70), .B(new_n206), .C1(new_n311), .C2(new_n313), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n304), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT71), .B1(new_n267), .B2(new_n281), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n279), .A2(new_n280), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n294), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n323), .A2(new_n326), .A3(KEYINPUT30), .A4(new_n291), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n298), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n316), .A2(new_n321), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n326), .A3(new_n329), .A4(new_n291), .ZN(new_n330));
  INV_X1    g144(.A(G237), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n188), .A3(G210), .ZN(new_n332));
  INV_X1    g146(.A(G101), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n334), .B(new_n335), .Z(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT31), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n328), .A2(KEYINPUT31), .A3(new_n330), .A4(new_n336), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n329), .B(new_n291), .C1(new_n281), .C2(new_n267), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n296), .A2(new_n322), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(new_n330), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n343), .ZN(new_n347));
  INV_X1    g161(.A(new_n336), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(G472), .A2(G902), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT32), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n339), .A2(new_n340), .B1(new_n347), .B2(new_n348), .ZN(new_n354));
  INV_X1    g168(.A(new_n351), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n356), .A3(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n350), .A2(new_n351), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n353), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n328), .A2(new_n330), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n348), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(new_n347), .C2(new_n348), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n323), .A2(new_n326), .A3(new_n291), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n322), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n330), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT28), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n344), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n336), .A2(KEYINPUT29), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT73), .B(new_n231), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n343), .B1(new_n367), .B2(new_n330), .ZN(new_n374));
  INV_X1    g188(.A(new_n344), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(new_n371), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n373), .B1(new_n376), .B2(G902), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n365), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n378), .A2(G472), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n245), .B1(new_n361), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n188), .A2(G227), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G101), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n386), .A2(new_n389), .A3(new_n333), .A4(new_n390), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n294), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n208), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n284), .B1(new_n259), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n390), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n385), .A2(G107), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n395), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n287), .A2(KEYINPUT10), .A3(new_n404), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n397), .A2(new_n281), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n403), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n411), .A2(KEYINPUT12), .A3(new_n324), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT12), .B1(new_n411), .B2(new_n324), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n384), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT81), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n409), .A2(new_n384), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n397), .A2(new_n407), .A3(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n324), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n409), .A2(KEYINPUT82), .A3(new_n384), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(G469), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G469), .A2(G902), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n412), .A2(new_n413), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n419), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n384), .B1(new_n423), .B2(new_n409), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n428), .B(new_n231), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT9), .B(G234), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G221), .B1(new_n435), .B2(G902), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n385), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n331), .A2(new_n188), .A3(G214), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n250), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n331), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(KEYINPUT18), .A2(G131), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT89), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(KEYINPUT18), .A3(G131), .ZN(new_n452));
  OR3_X1    g266(.A1(new_n200), .A2(KEYINPUT88), .A3(new_n202), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT88), .B1(new_n200), .B2(new_n202), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n224), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n445), .A2(new_n277), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n444), .A2(new_n458), .A3(G131), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n444), .B2(G131), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n193), .A3(new_n223), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT19), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(new_n200), .ZN(new_n466));
  INV_X1    g280(.A(new_n222), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n462), .A2(new_n468), .A3(new_n221), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n440), .B1(new_n456), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n461), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT17), .A3(new_n459), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n203), .B(new_n472), .C1(new_n462), .C2(KEYINPUT17), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n439), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n231), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT20), .ZN(new_n479));
  AOI21_X1  g293(.A(G475), .B1(new_n470), .B2(new_n475), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n231), .ZN(new_n482));
  INV_X1    g296(.A(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n439), .B1(new_n473), .B2(new_n474), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n231), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n479), .A2(new_n482), .B1(G475), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n188), .A2(G952), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(G234), .B2(G237), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT21), .B(G898), .Z(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n231), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n494));
  INV_X1    g308(.A(G122), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n308), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n310), .A2(G122), .ZN(new_n497));
  OR3_X1    g311(.A1(new_n496), .A2(KEYINPUT14), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(KEYINPUT14), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(G107), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n496), .A2(new_n497), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n388), .ZN(new_n502));
  XNOR2_X1  g316(.A(G128), .B(G143), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n269), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(KEYINPUT13), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n208), .A2(KEYINPUT13), .A3(G143), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n269), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n506), .A2(new_n508), .B1(new_n269), .B2(new_n503), .ZN(new_n509));
  INV_X1    g323(.A(new_n502), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n501), .A2(new_n388), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n435), .A2(new_n230), .A3(G953), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n505), .B2(new_n512), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n494), .B(new_n231), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n505), .A2(new_n512), .ZN(new_n521));
  INV_X1    g335(.A(new_n513), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  INV_X1    g338(.A(new_n519), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n494), .A3(new_n231), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n487), .A2(new_n493), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT5), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n309), .B2(new_n315), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n531));
  OAI21_X1  g345(.A(G113), .B1(new_n531), .B2(new_n317), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n321), .B(new_n404), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT5), .B1(new_n319), .B2(new_n320), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT86), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n321), .A4(new_n404), .ZN(new_n539));
  INV_X1    g353(.A(new_n531), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n309), .B2(new_n315), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n321), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n403), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(G110), .B(G122), .Z(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n396), .A2(new_n393), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT83), .B1(new_n329), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n322), .A2(new_n550), .A3(new_n393), .A4(new_n396), .ZN(new_n551));
  INV_X1    g365(.A(new_n545), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n321), .B(new_n404), .C1(new_n541), .C2(new_n532), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n549), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT85), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n294), .B2(new_n198), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n267), .A2(KEYINPUT85), .A3(G125), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n198), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n558));
  INV_X1    g372(.A(G224), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G953), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n294), .B2(new_n198), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n561), .B2(new_n560), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n547), .A2(new_n554), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n231), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n553), .A3(new_n551), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n545), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT6), .A3(new_n554), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n560), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT6), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n575), .A3(new_n545), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n566), .A2(KEYINPUT87), .A3(new_n231), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G210), .B1(G237), .B2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n569), .A2(new_n577), .A3(new_n580), .A4(new_n578), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G214), .B1(G237), .B2(G902), .ZN(new_n585));
  AND4_X1   g399(.A1(new_n437), .A2(new_n528), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n381), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT93), .B(G101), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G3));
  INV_X1    g403(.A(new_n585), .ZN(new_n590));
  AND4_X1   g404(.A1(new_n580), .A2(new_n569), .A3(new_n577), .A4(new_n578), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(KEYINPUT94), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n582), .A2(new_n593), .A3(new_n583), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n592), .A2(KEYINPUT95), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT95), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(new_n596), .A3(new_n493), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n524), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT33), .B1(new_n523), .B2(new_n514), .ZN(new_n600));
  OAI21_X1  g414(.A(G478), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n524), .A2(new_n518), .A3(new_n231), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n518), .A2(new_n231), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n486), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G472), .B1(new_n354), .B2(G902), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n437), .A2(new_n608), .A3(new_n358), .A4(new_n244), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT34), .B(G104), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(new_n609), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n485), .A2(G475), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n480), .A2(new_n481), .A3(new_n231), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n481), .B1(new_n480), .B2(new_n231), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n527), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n597), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT96), .Z(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  AND2_X1   g436(.A1(new_n608), .A2(new_n358), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n227), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n234), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n243), .A2(new_n233), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n586), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G12));
  INV_X1    g447(.A(new_n437), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n361), .B2(new_n380), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n595), .A2(new_n596), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n489), .B1(new_n492), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n635), .A2(new_n636), .A3(new_n630), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  INV_X1    g455(.A(G472), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n362), .A2(new_n336), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n231), .B1(new_n368), .B2(new_n336), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n642), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n361), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n630), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n486), .B1(new_n520), .B2(new_n526), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n585), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n584), .B(KEYINPUT38), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n649), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT98), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n638), .B(KEYINPUT39), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n634), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G143), .ZN(G45));
  INV_X1    g473(.A(new_n638), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n606), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n635), .A2(new_n636), .A3(new_n630), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  OR2_X1    g478(.A1(new_n430), .A2(new_n431), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n231), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G469), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n432), .ZN(new_n668));
  INV_X1    g482(.A(new_n436), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n597), .A2(new_n381), .A3(new_n606), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  INV_X1    g487(.A(new_n670), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n595), .A2(new_n596), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n361), .A2(new_n380), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n493), .B(new_n236), .C1(new_n243), .C2(new_n233), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n618), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND4_X1  g493(.A1(new_n675), .A2(new_n676), .A3(new_n528), .A4(new_n630), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n369), .A2(new_n682), .A3(new_n344), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT99), .B1(new_n374), .B2(new_n375), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n348), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n341), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT100), .B1(new_n686), .B2(new_n351), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  AOI211_X1 g502(.A(new_n688), .B(new_n355), .C1(new_n341), .C2(new_n685), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n677), .B(new_n608), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n636), .A2(new_n691), .A3(new_n650), .A4(new_n670), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G122), .ZN(G24));
  OAI211_X1 g507(.A(new_n608), .B(new_n630), .C1(new_n687), .C2(new_n689), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n662), .B(new_n675), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n379), .B1(new_n357), .B2(new_n360), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n582), .A2(new_n583), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n427), .B(KEYINPUT102), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n425), .A2(KEYINPUT103), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n425), .A2(KEYINPUT103), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n418), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n432), .B(new_n703), .C1(new_n706), .C2(new_n428), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n669), .A2(new_n590), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n701), .A2(new_n245), .A3(new_n661), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n700), .B1(new_n710), .B2(KEYINPUT42), .ZN(new_n711));
  INV_X1    g525(.A(new_n709), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n381), .A2(new_n662), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(KEYINPUT104), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n709), .A2(new_n661), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n380), .A2(new_n356), .A3(new_n352), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n244), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G131), .ZN(G33));
  AND3_X1   g535(.A1(new_n381), .A2(new_n639), .A3(new_n712), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n269), .ZN(G36));
  OAI211_X1 g537(.A(KEYINPUT45), .B(new_n418), .C1(new_n704), .C2(new_n705), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT45), .B1(new_n418), .B2(new_n425), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n428), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n703), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n432), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT46), .B1(new_n729), .B2(new_n703), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n436), .ZN(new_n734));
  INV_X1    g548(.A(new_n605), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n486), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n736), .B1(KEYINPUT106), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n623), .B1(new_n742), .B2(KEYINPUT107), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n741), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n649), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT44), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n734), .A2(new_n655), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n743), .A2(KEYINPUT44), .A3(new_n746), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n584), .A2(new_n590), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT108), .Z(new_n751));
  AOI21_X1  g565(.A(KEYINPUT109), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n751), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n748), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n734), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n436), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n661), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n676), .A2(new_n244), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT110), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n761), .A2(new_n765), .A3(new_n750), .A4(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NOR3_X1   g582(.A1(new_n649), .A2(new_n527), .A3(new_n487), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n635), .A2(new_n660), .A3(new_n750), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT113), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n701), .A2(new_n634), .A3(new_n638), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n750), .A4(new_n769), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n617), .B1(new_n486), .B2(new_n605), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n584), .A2(new_n776), .A3(new_n585), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n609), .A2(new_n777), .A3(new_n493), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n381), .B2(new_n586), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n678), .A2(new_n680), .A3(new_n779), .A4(new_n692), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n671), .A2(new_n631), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n775), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n696), .A2(new_n697), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n717), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n722), .B1(new_n716), .B2(new_n719), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n698), .A2(new_n640), .A3(new_n663), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n648), .A2(new_n436), .A3(new_n649), .A4(new_n660), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n592), .A2(new_n594), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n592), .A2(new_n594), .A3(KEYINPUT95), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n650), .A4(new_n707), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n788), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n646), .B1(new_n357), .B2(new_n360), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n630), .A3(new_n638), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n792), .A2(new_n793), .A3(new_n650), .A4(new_n707), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT114), .A4(new_n436), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(new_n787), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n787), .A2(new_n800), .A3(KEYINPUT52), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n787), .A2(new_n800), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n786), .B(KEYINPUT53), .C1(new_n804), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n787), .A2(new_n800), .A3(KEYINPUT52), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n801), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n782), .A2(new_n785), .A3(new_n784), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n805), .A2(new_n806), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n812), .B2(KEYINPUT115), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n814), .B1(new_n818), .B2(new_n807), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(KEYINPUT117), .A3(KEYINPUT53), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n813), .A2(new_n814), .A3(new_n811), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n786), .B1(new_n804), .B2(new_n808), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n811), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n824), .B1(new_n827), .B2(new_n822), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n819), .A2(KEYINPUT53), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n829), .C2(new_n825), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n744), .A2(new_n489), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n608), .B1(new_n687), .B2(new_n689), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n245), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n670), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n652), .A2(new_n585), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n835), .A2(KEYINPUT50), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n750), .A2(new_n489), .A3(new_n670), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n742), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n783), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT50), .B1(new_n835), .B2(new_n837), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n648), .A2(new_n245), .A3(new_n839), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n486), .A3(new_n605), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n841), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n667), .A2(new_n669), .A3(new_n432), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n759), .A2(new_n760), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n834), .A2(new_n751), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n847), .A2(new_n852), .B1(new_n606), .B2(new_n844), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n759), .A2(new_n760), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n759), .A2(new_n856), .A3(new_n760), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n849), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n846), .B1(new_n858), .B2(new_n851), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n853), .B1(new_n859), .B2(KEYINPUT51), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n675), .B2(new_n834), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n840), .A2(new_n244), .A3(new_n718), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT48), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n488), .B(KEYINPUT119), .Z(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n831), .A2(new_n865), .B1(G952), .B2(G953), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n668), .A2(KEYINPUT49), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n737), .A2(new_n867), .A3(new_n244), .A4(new_n708), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n652), .B1(new_n868), .B2(KEYINPUT111), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(KEYINPUT111), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n668), .A2(KEYINPUT49), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT112), .Z(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n796), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n188), .A2(G952), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT120), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n816), .A2(new_n820), .A3(G210), .A4(G902), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n572), .A2(new_n576), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n574), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n882), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n876), .B1(new_n883), .B2(new_n884), .ZN(G51));
  XOR2_X1   g699(.A(new_n703), .B(KEYINPUT57), .Z(new_n886));
  AND3_X1   g700(.A1(new_n816), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT54), .B1(new_n816), .B2(new_n820), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n665), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n821), .A2(new_n231), .A3(new_n729), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n875), .B1(new_n890), .B2(new_n891), .ZN(G54));
  INV_X1    g706(.A(new_n875), .ZN(new_n893));
  AND2_X1   g707(.A1(KEYINPUT58), .A2(G475), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n816), .A2(new_n820), .A3(G902), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n476), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n898), .A2(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(KEYINPUT121), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(G60));
  NOR2_X1   g715(.A1(new_n599), .A2(new_n600), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n604), .B(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n831), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n902), .B(new_n904), .C1(new_n887), .C2(new_n888), .ZN(new_n906));
  INV_X1    g720(.A(new_n876), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n908), .ZN(G63));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n230), .A2(new_n231), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n816), .A2(new_n820), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n229), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n627), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n907), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n910), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n914), .A2(new_n917), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(KEYINPUT61), .A3(new_n907), .A4(new_n915), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G66));
  OAI21_X1  g736(.A(G953), .B1(new_n491), .B2(new_n559), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n780), .A2(new_n781), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n880), .B1(G898), .B2(new_n188), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  AOI21_X1  g741(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n718), .A2(new_n244), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n734), .A2(new_n655), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n636), .A3(new_n650), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n756), .A2(new_n931), .A3(new_n787), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n764), .B2(new_n766), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n785), .B(KEYINPUT125), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n188), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n298), .A2(new_n327), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n466), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n935), .B(new_n937), .C1(new_n637), .C2(new_n188), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n928), .B1(new_n938), .B2(KEYINPUT124), .ZN(new_n939));
  INV_X1    g753(.A(new_n937), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n658), .A2(new_n787), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n658), .A2(KEYINPUT62), .A3(new_n787), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n945), .A2(new_n756), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n381), .A2(new_n656), .A3(new_n750), .A4(new_n776), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n764), .B2(new_n766), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n940), .B1(new_n950), .B2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n938), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n939), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n951), .B(new_n938), .C1(KEYINPUT124), .C2(new_n928), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G72));
  NAND3_X1  g769(.A1(new_n946), .A2(new_n949), .A3(new_n924), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n642), .A2(new_n231), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n643), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n956), .A2(KEYINPUT127), .A3(new_n959), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n363), .A2(new_n337), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n959), .C1(new_n829), .C2(new_n825), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n933), .A2(new_n924), .A3(new_n934), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n336), .B1(new_n968), .B2(new_n959), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n330), .A3(new_n328), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n893), .A2(new_n965), .A3(new_n967), .A4(new_n970), .ZN(G57));
endmodule


