

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752;

  XNOR2_X2 U375 ( .A(n435), .B(n717), .ZN(n451) );
  XNOR2_X2 U376 ( .A(n366), .B(n421), .ZN(n435) );
  NOR2_X2 U377 ( .A1(n365), .A2(n561), .ZN(n440) );
  OR2_X1 U378 ( .A1(n619), .A2(n525), .ZN(n390) );
  XNOR2_X1 U379 ( .A(n511), .B(n510), .ZN(n619) );
  OR2_X1 U380 ( .A1(n515), .A2(n502), .ZN(n504) );
  AND2_X1 U381 ( .A1(n395), .A2(n394), .ZN(n393) );
  OR2_X1 U382 ( .A1(n676), .A2(n392), .ZN(n391) );
  XNOR2_X1 U383 ( .A(n420), .B(n419), .ZN(n627) );
  XNOR2_X1 U384 ( .A(n737), .B(G101), .ZN(n366) );
  XNOR2_X1 U385 ( .A(G116), .B(KEYINPUT3), .ZN(n384) );
  INV_X2 U386 ( .A(KEYINPUT4), .ZN(n367) );
  INV_X2 U387 ( .A(G953), .ZN(n725) );
  AND2_X1 U388 ( .A1(n354), .A2(n355), .ZN(n529) );
  NAND2_X1 U389 ( .A1(n512), .A2(n358), .ZN(n354) );
  XOR2_X1 U390 ( .A(n385), .B(KEYINPUT100), .Z(n355) );
  NOR2_X1 U391 ( .A1(n616), .A2(n716), .ZN(n618) );
  NAND2_X1 U392 ( .A1(n505), .A2(n629), .ZN(n365) );
  AND2_X2 U393 ( .A1(n620), .A2(n605), .ZN(n357) );
  NOR2_X2 U394 ( .A1(G902), .A2(n707), .ZN(n428) );
  XNOR2_X2 U395 ( .A(n518), .B(KEYINPUT1), .ZN(n505) );
  XNOR2_X2 U396 ( .A(n428), .B(n427), .ZN(n518) );
  XNOR2_X1 U397 ( .A(n382), .B(n585), .ZN(n586) );
  XNOR2_X1 U398 ( .A(n447), .B(n404), .ZN(n472) );
  BUF_X1 U399 ( .A(n518), .Z(n544) );
  NOR2_X1 U400 ( .A1(n626), .A2(n627), .ZN(n629) );
  NAND2_X1 U401 ( .A1(n356), .A2(n388), .ZN(n387) );
  INV_X1 U402 ( .A(n573), .ZN(n388) );
  XNOR2_X1 U403 ( .A(n403), .B(G125), .ZN(n447) );
  NOR2_X1 U404 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U405 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U406 ( .A(n738), .ZN(n376) );
  XNOR2_X1 U407 ( .A(n470), .B(n469), .ZN(n515) );
  XNOR2_X1 U408 ( .A(n380), .B(KEYINPUT39), .ZN(n598) );
  NAND2_X1 U409 ( .A1(n378), .A2(n550), .ZN(n380) );
  NOR2_X1 U410 ( .A1(n552), .A2(n379), .ZN(n378) );
  XNOR2_X1 U411 ( .A(n487), .B(n486), .ZN(n514) );
  XNOR2_X1 U412 ( .A(n485), .B(KEYINPUT13), .ZN(n486) );
  INV_X1 U413 ( .A(G475), .ZN(n485) );
  NAND2_X1 U414 ( .A1(n371), .A2(KEYINPUT70), .ZN(n370) );
  INV_X1 U415 ( .A(n749), .ZN(n372) );
  NAND2_X1 U416 ( .A1(n390), .A2(KEYINPUT64), .ZN(n389) );
  NAND2_X1 U417 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U418 ( .A(G469), .ZN(n427) );
  OR2_X1 U419 ( .A1(n603), .A2(n599), .ZN(n738) );
  XNOR2_X1 U420 ( .A(G119), .B(G128), .ZN(n408) );
  INV_X1 U421 ( .A(KEYINPUT89), .ZN(n406) );
  XNOR2_X1 U422 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n405) );
  XNOR2_X1 U423 ( .A(n446), .B(G134), .ZN(n494) );
  NAND2_X1 U424 ( .A1(n374), .A2(n373), .ZN(n606) );
  INV_X1 U425 ( .A(KEYINPUT2), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n582), .B(n581), .ZN(n639) );
  XNOR2_X1 U427 ( .A(n579), .B(n383), .ZN(n747) );
  XNOR2_X1 U428 ( .A(n521), .B(KEYINPUT93), .ZN(n686) );
  NAND2_X1 U429 ( .A1(n360), .A2(n393), .ZN(n566) );
  OR2_X1 U430 ( .A1(n698), .A2(n686), .ZN(n356) );
  XNOR2_X1 U431 ( .A(n566), .B(KEYINPUT19), .ZN(n546) );
  AND2_X1 U432 ( .A1(n369), .A2(n368), .ZN(n358) );
  XNOR2_X1 U433 ( .A(n531), .B(n530), .ZN(n724) );
  INV_X1 U434 ( .A(n724), .ZN(n375) );
  XNOR2_X1 U435 ( .A(G143), .B(G128), .ZN(n446) );
  AND2_X1 U436 ( .A1(n749), .A2(KEYINPUT44), .ZN(n359) );
  AND2_X1 U437 ( .A1(n391), .A2(n643), .ZN(n360) );
  XOR2_X1 U438 ( .A(n608), .B(n607), .Z(n361) );
  AND2_X1 U439 ( .A1(KEYINPUT64), .A2(KEYINPUT70), .ZN(n362) );
  AND2_X1 U440 ( .A1(n370), .A2(KEYINPUT64), .ZN(n363) );
  XOR2_X1 U441 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n364) );
  NOR2_X1 U442 ( .A1(n365), .A2(n542), .ZN(n637) );
  XNOR2_X2 U443 ( .A(n367), .B(KEYINPUT71), .ZN(n737) );
  NAND2_X1 U444 ( .A1(n749), .A2(n363), .ZN(n368) );
  NAND2_X1 U445 ( .A1(n372), .A2(n362), .ZN(n369) );
  INV_X1 U446 ( .A(KEYINPUT44), .ZN(n371) );
  NAND2_X1 U447 ( .A1(n374), .A2(n364), .ZN(n621) );
  AND2_X1 U448 ( .A1(n377), .A2(n550), .ZN(n577) );
  NOR2_X1 U449 ( .A1(n552), .A2(n381), .ZN(n377) );
  NAND2_X1 U450 ( .A1(n644), .A2(n551), .ZN(n379) );
  INV_X1 U451 ( .A(n551), .ZN(n381) );
  NAND2_X1 U452 ( .A1(n751), .A2(n747), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n578), .B(KEYINPUT107), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(G119), .ZN(n431) );
  INV_X1 U455 ( .A(n684), .ZN(n386) );
  NAND2_X1 U456 ( .A1(n389), .A2(n359), .ZN(n527) );
  NAND2_X1 U457 ( .A1(n393), .A2(n391), .ZN(n595) );
  OR2_X1 U458 ( .A1(n458), .A2(n605), .ZN(n392) );
  NAND2_X1 U459 ( .A1(n458), .A2(n605), .ZN(n394) );
  NAND2_X1 U460 ( .A1(n676), .A2(n458), .ZN(n395) );
  BUF_X1 U461 ( .A(n705), .Z(n711) );
  AND2_X2 U462 ( .A1(n606), .A2(n357), .ZN(n705) );
  NAND2_X1 U463 ( .A1(n705), .A2(G472), .ZN(n609) );
  OR2_X1 U464 ( .A1(G902), .A2(n614), .ZN(n396) );
  XOR2_X1 U465 ( .A(n407), .B(n406), .Z(n397) );
  AND2_X1 U466 ( .A1(n627), .A2(n505), .ZN(n398) );
  INV_X1 U467 ( .A(n639), .ZN(n640) );
  NOR2_X1 U468 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U469 ( .A(KEYINPUT10), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n397), .B(n410), .ZN(n411) );
  NOR2_X1 U471 ( .A1(n565), .A2(n564), .ZN(n590) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n419) );
  INV_X1 U473 ( .A(n716), .ZN(n611) );
  XNOR2_X1 U474 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U475 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U476 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n400) );
  XNOR2_X1 U477 ( .A(G902), .B(KEYINPUT15), .ZN(n453) );
  NAND2_X1 U478 ( .A1(G234), .A2(n453), .ZN(n399) );
  XNOR2_X1 U479 ( .A(n400), .B(n399), .ZN(n416) );
  AND2_X1 U480 ( .A1(n416), .A2(G221), .ZN(n402) );
  INV_X1 U481 ( .A(KEYINPUT21), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n402), .B(n401), .ZN(n626) );
  INV_X1 U483 ( .A(G146), .ZN(n403) );
  XNOR2_X1 U484 ( .A(n472), .B(n405), .ZN(n412) );
  XNOR2_X1 U485 ( .A(G110), .B(G137), .ZN(n407) );
  XOR2_X1 U486 ( .A(KEYINPUT90), .B(G140), .Z(n409) );
  XNOR2_X1 U487 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U488 ( .A(n412), .B(n411), .ZN(n415) );
  NAND2_X1 U489 ( .A1(G234), .A2(n725), .ZN(n413) );
  XOR2_X1 U490 ( .A(KEYINPUT8), .B(n413), .Z(n495) );
  NAND2_X1 U491 ( .A1(G221), .A2(n495), .ZN(n414) );
  XNOR2_X1 U492 ( .A(n415), .B(n414), .ZN(n712) );
  NOR2_X1 U493 ( .A1(G902), .A2(n712), .ZN(n420) );
  AND2_X1 U494 ( .A1(G217), .A2(n416), .ZN(n418) );
  XNOR2_X1 U495 ( .A(KEYINPUT25), .B(KEYINPUT92), .ZN(n417) );
  XOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n421) );
  XOR2_X1 U497 ( .A(G104), .B(G110), .Z(n422) );
  XNOR2_X1 U498 ( .A(n422), .B(G107), .ZN(n717) );
  XOR2_X1 U499 ( .A(G140), .B(G131), .Z(n473) );
  XOR2_X1 U500 ( .A(n473), .B(KEYINPUT74), .Z(n424) );
  NAND2_X1 U501 ( .A1(G227), .A2(n725), .ZN(n423) );
  XNOR2_X1 U502 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U503 ( .A(n451), .B(n425), .ZN(n426) );
  XNOR2_X1 U504 ( .A(n494), .B(G137), .ZN(n734) );
  XNOR2_X1 U505 ( .A(G146), .B(n734), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n426), .B(n438), .ZN(n707) );
  INV_X1 U507 ( .A(KEYINPUT73), .ZN(n429) );
  XNOR2_X1 U508 ( .A(n429), .B(G113), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n431), .B(n430), .ZN(n442) );
  XOR2_X1 U510 ( .A(G131), .B(KEYINPUT5), .Z(n433) );
  NOR2_X1 U511 ( .A1(G953), .A2(G237), .ZN(n474) );
  NAND2_X1 U512 ( .A1(n474), .A2(G210), .ZN(n432) );
  XNOR2_X1 U513 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U514 ( .A(n442), .B(n434), .ZN(n436) );
  XNOR2_X1 U515 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U516 ( .A(n438), .B(n437), .ZN(n608) );
  INV_X1 U517 ( .A(G902), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n608), .A2(n455), .ZN(n439) );
  XNOR2_X2 U519 ( .A(n439), .B(G472), .ZN(n635) );
  XNOR2_X1 U520 ( .A(n635), .B(KEYINPUT6), .ZN(n561) );
  XNOR2_X1 U521 ( .A(n440), .B(KEYINPUT33), .ZN(n622) );
  XNOR2_X1 U522 ( .A(KEYINPUT16), .B(G122), .ZN(n441) );
  XNOR2_X1 U523 ( .A(n442), .B(n441), .ZN(n718) );
  XOR2_X1 U524 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n445) );
  NAND2_X1 U525 ( .A1(G224), .A2(n725), .ZN(n443) );
  XNOR2_X1 U526 ( .A(n443), .B(KEYINPUT75), .ZN(n444) );
  XNOR2_X1 U527 ( .A(n445), .B(n444), .ZN(n449) );
  XNOR2_X1 U528 ( .A(n446), .B(n447), .ZN(n448) );
  XNOR2_X1 U529 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U530 ( .A(n718), .B(n450), .ZN(n452) );
  XNOR2_X1 U531 ( .A(n452), .B(n451), .ZN(n676) );
  INV_X1 U532 ( .A(n453), .ZN(n605) );
  INV_X1 U533 ( .A(G237), .ZN(n454) );
  NAND2_X1 U534 ( .A1(n455), .A2(n454), .ZN(n459) );
  NAND2_X1 U535 ( .A1(n459), .A2(G210), .ZN(n457) );
  XNOR2_X1 U536 ( .A(KEYINPUT77), .B(KEYINPUT87), .ZN(n456) );
  XNOR2_X1 U537 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U538 ( .A1(n459), .A2(G214), .ZN(n643) );
  NAND2_X1 U539 ( .A1(G234), .A2(G237), .ZN(n460) );
  XNOR2_X1 U540 ( .A(n460), .B(KEYINPUT14), .ZN(n463) );
  NAND2_X1 U541 ( .A1(G952), .A2(n463), .ZN(n461) );
  XOR2_X1 U542 ( .A(KEYINPUT88), .B(n461), .Z(n660) );
  NAND2_X1 U543 ( .A1(n660), .A2(n725), .ZN(n532) );
  AND2_X1 U544 ( .A1(G953), .A2(G902), .ZN(n462) );
  NAND2_X1 U545 ( .A1(n463), .A2(n462), .ZN(n533) );
  INV_X1 U546 ( .A(n533), .ZN(n465) );
  INV_X1 U547 ( .A(G898), .ZN(n464) );
  NAND2_X1 U548 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U549 ( .A1(n532), .A2(n466), .ZN(n467) );
  NAND2_X1 U550 ( .A1(n546), .A2(n467), .ZN(n470) );
  INV_X1 U551 ( .A(KEYINPUT67), .ZN(n468) );
  XNOR2_X1 U552 ( .A(n468), .B(KEYINPUT0), .ZN(n469) );
  NOR2_X1 U553 ( .A1(n622), .A2(n515), .ZN(n471) );
  XNOR2_X1 U554 ( .A(n471), .B(KEYINPUT34), .ZN(n498) );
  XOR2_X1 U555 ( .A(n473), .B(n472), .Z(n733) );
  XOR2_X1 U556 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n476) );
  NAND2_X1 U557 ( .A1(n474), .A2(G214), .ZN(n475) );
  XNOR2_X1 U558 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U559 ( .A(n477), .B(KEYINPUT97), .Z(n483) );
  XOR2_X1 U560 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n479) );
  XNOR2_X1 U561 ( .A(G122), .B(G143), .ZN(n478) );
  XNOR2_X1 U562 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U563 ( .A(G104), .B(G113), .ZN(n480) );
  XNOR2_X1 U564 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U565 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U566 ( .A(n733), .B(n484), .ZN(n671) );
  NOR2_X1 U567 ( .A1(G902), .A2(n671), .ZN(n487) );
  XOR2_X1 U568 ( .A(KEYINPUT99), .B(KEYINPUT7), .Z(n489) );
  XNOR2_X1 U569 ( .A(G122), .B(KEYINPUT9), .ZN(n488) );
  XNOR2_X1 U570 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U571 ( .A(n490), .B(KEYINPUT98), .Z(n492) );
  XNOR2_X1 U572 ( .A(G107), .B(G116), .ZN(n491) );
  XNOR2_X1 U573 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U574 ( .A(n494), .B(n493), .Z(n497) );
  NAND2_X1 U575 ( .A1(G217), .A2(n495), .ZN(n496) );
  XNOR2_X1 U576 ( .A(n497), .B(n496), .ZN(n614) );
  XNOR2_X1 U577 ( .A(G478), .B(n396), .ZN(n513) );
  INV_X1 U578 ( .A(n513), .ZN(n501) );
  NOR2_X1 U579 ( .A1(n514), .A2(n501), .ZN(n553) );
  NAND2_X1 U580 ( .A1(n498), .A2(n553), .ZN(n500) );
  XOR2_X1 U581 ( .A(KEYINPUT76), .B(KEYINPUT35), .Z(n499) );
  XNOR2_X2 U582 ( .A(n500), .B(n499), .ZN(n749) );
  AND2_X1 U583 ( .A1(n514), .A2(n501), .ZN(n580) );
  INV_X1 U584 ( .A(n626), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n580), .A2(n537), .ZN(n502) );
  INV_X1 U586 ( .A(KEYINPUT22), .ZN(n503) );
  XNOR2_X2 U587 ( .A(n504), .B(n503), .ZN(n508) );
  NOR2_X1 U588 ( .A1(n505), .A2(n635), .ZN(n506) );
  AND2_X1 U589 ( .A1(n627), .A2(n506), .ZN(n507) );
  AND2_X1 U590 ( .A1(n508), .A2(n507), .ZN(n690) );
  NAND2_X1 U591 ( .A1(n508), .A2(n561), .ZN(n523) );
  INV_X1 U592 ( .A(n523), .ZN(n509) );
  NAND2_X1 U593 ( .A1(n509), .A2(n398), .ZN(n511) );
  XNOR2_X1 U594 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n510) );
  NOR2_X1 U595 ( .A1(n690), .A2(n619), .ZN(n512) );
  NOR2_X1 U596 ( .A1(n514), .A2(n513), .ZN(n696) );
  AND2_X1 U597 ( .A1(n514), .A2(n513), .ZN(n699) );
  NOR2_X1 U598 ( .A1(n696), .A2(n699), .ZN(n648) );
  XOR2_X1 U599 ( .A(n648), .B(KEYINPUT83), .Z(n573) );
  XOR2_X1 U600 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n517) );
  INV_X1 U601 ( .A(n635), .ZN(n542) );
  INV_X1 U602 ( .A(n515), .ZN(n519) );
  NAND2_X1 U603 ( .A1(n637), .A2(n519), .ZN(n516) );
  XOR2_X1 U604 ( .A(n517), .B(n516), .Z(n698) );
  NAND2_X1 U605 ( .A1(n544), .A2(n629), .ZN(n552) );
  NOR2_X1 U606 ( .A1(n552), .A2(n635), .ZN(n520) );
  NAND2_X1 U607 ( .A1(n520), .A2(n519), .ZN(n521) );
  INV_X1 U608 ( .A(n627), .ZN(n539) );
  INV_X1 U609 ( .A(n505), .ZN(n570) );
  NAND2_X1 U610 ( .A1(n539), .A2(n570), .ZN(n522) );
  NOR2_X1 U611 ( .A1(n523), .A2(n522), .ZN(n684) );
  INV_X1 U612 ( .A(n690), .ZN(n524) );
  NAND2_X1 U613 ( .A1(n524), .A2(KEYINPUT70), .ZN(n525) );
  NAND2_X1 U614 ( .A1(n371), .A2(KEYINPUT64), .ZN(n526) );
  NAND2_X1 U615 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n529), .A2(n528), .ZN(n531) );
  XOR2_X1 U617 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n530) );
  INV_X1 U618 ( .A(n532), .ZN(n656) );
  XOR2_X1 U619 ( .A(n533), .B(KEYINPUT101), .Z(n534) );
  NOR2_X1 U620 ( .A1(G900), .A2(n534), .ZN(n535) );
  NOR2_X1 U621 ( .A1(n656), .A2(n535), .ZN(n536) );
  XOR2_X1 U622 ( .A(KEYINPUT78), .B(n536), .Z(n551) );
  NAND2_X1 U623 ( .A1(n537), .A2(n551), .ZN(n538) );
  INV_X1 U624 ( .A(KEYINPUT72), .ZN(n540) );
  XNOR2_X1 U625 ( .A(n541), .B(n540), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n562), .A2(n542), .ZN(n543) );
  XNOR2_X1 U627 ( .A(n543), .B(KEYINPUT28), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n583) );
  INV_X1 U629 ( .A(n583), .ZN(n547) );
  NAND2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n572), .A2(KEYINPUT47), .ZN(n548) );
  XNOR2_X1 U632 ( .A(n548), .B(KEYINPUT82), .ZN(n559) );
  AND2_X1 U633 ( .A1(n648), .A2(KEYINPUT47), .ZN(n557) );
  NAND2_X1 U634 ( .A1(n635), .A2(n643), .ZN(n549) );
  XOR2_X1 U635 ( .A(KEYINPUT30), .B(n549), .Z(n550) );
  INV_X1 U636 ( .A(n553), .ZN(n554) );
  NOR2_X1 U637 ( .A1(n554), .A2(n595), .ZN(n555) );
  NAND2_X1 U638 ( .A1(n577), .A2(n555), .ZN(n556) );
  XNOR2_X1 U639 ( .A(KEYINPUT105), .B(n556), .ZN(n748) );
  NOR2_X1 U640 ( .A1(n557), .A2(n748), .ZN(n558) );
  AND2_X1 U641 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U642 ( .A(n560), .B(KEYINPUT81), .ZN(n571) );
  INV_X1 U643 ( .A(n696), .ZN(n565) );
  OR2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U645 ( .A(KEYINPUT102), .B(n563), .ZN(n564) );
  INV_X1 U646 ( .A(n566), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n590), .A2(n567), .ZN(n568) );
  XNOR2_X1 U648 ( .A(n568), .B(KEYINPUT36), .ZN(n569) );
  NOR2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n702) );
  NOR2_X1 U650 ( .A1(n571), .A2(n702), .ZN(n576) );
  INV_X1 U651 ( .A(n572), .ZN(n693) );
  NOR2_X1 U652 ( .A1(KEYINPUT47), .A2(n573), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n693), .A2(n574), .ZN(n575) );
  NAND2_X1 U654 ( .A1(n576), .A2(n575), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n595), .B(KEYINPUT38), .ZN(n644) );
  NAND2_X1 U656 ( .A1(n696), .A2(n598), .ZN(n579) );
  XOR2_X1 U657 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n578) );
  NAND2_X1 U658 ( .A1(n644), .A2(n643), .ZN(n647) );
  INV_X1 U659 ( .A(n580), .ZN(n646) );
  NOR2_X1 U660 ( .A1(n647), .A2(n646), .ZN(n582) );
  XNOR2_X1 U661 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n581) );
  NOR2_X1 U662 ( .A1(n639), .A2(n583), .ZN(n584) );
  XOR2_X1 U663 ( .A(KEYINPUT42), .B(n584), .Z(n751) );
  XOR2_X1 U664 ( .A(KEYINPUT46), .B(KEYINPUT85), .Z(n585) );
  INV_X1 U665 ( .A(KEYINPUT48), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(n588), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n590), .A2(n643), .ZN(n591) );
  NOR2_X1 U668 ( .A1(n505), .A2(n591), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n593), .B(n592), .ZN(n594) );
  AND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U672 ( .A(KEYINPUT104), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n597), .B(n596), .ZN(n750) );
  NAND2_X1 U674 ( .A1(n598), .A2(n699), .ZN(n704) );
  NAND2_X1 U675 ( .A1(n750), .A2(n704), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n704), .A2(KEYINPUT2), .ZN(n600) );
  XNOR2_X1 U677 ( .A(n600), .B(KEYINPUT79), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n750), .A2(n601), .ZN(n602) );
  OR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X2 U680 ( .A1(n604), .A2(n724), .ZN(n620) );
  XNOR2_X1 U681 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n609), .B(n361), .ZN(n612) );
  INV_X1 U683 ( .A(G952), .ZN(n610) );
  AND2_X1 U684 ( .A1(n610), .A2(G953), .ZN(n716) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U687 ( .A1(n705), .A2(G478), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U689 ( .A(KEYINPUT119), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n618), .B(n617), .ZN(G63) );
  XOR2_X1 U691 ( .A(n619), .B(G119), .Z(G21) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n639), .A2(n622), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT115), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n665) );
  NAND2_X1 U696 ( .A1(n665), .A2(n725), .ZN(n658) );
  AND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U698 ( .A(KEYINPUT49), .B(n628), .ZN(n633) );
  OR2_X1 U699 ( .A1(n629), .A2(n505), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT50), .ZN(n631) );
  XNOR2_X1 U701 ( .A(KEYINPUT112), .B(n631), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U705 ( .A(n638), .B(KEYINPUT51), .ZN(n641) );
  NAND2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n642), .B(KEYINPUT113), .ZN(n654) );
  NOR2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U709 ( .A1(n646), .A2(n645), .ZN(n651) );
  NOR2_X1 U710 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U711 ( .A(n649), .B(KEYINPUT114), .ZN(n650) );
  NOR2_X1 U712 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U713 ( .A1(n622), .A2(n652), .ZN(n653) );
  NOR2_X1 U714 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U715 ( .A(KEYINPUT52), .B(n655), .Z(n661) );
  NAND2_X1 U716 ( .A1(n661), .A2(n656), .ZN(n657) );
  AND2_X1 U717 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U718 ( .A1(n659), .A2(KEYINPUT116), .ZN(n667) );
  NAND2_X1 U719 ( .A1(n661), .A2(n660), .ZN(n663) );
  AND2_X1 U720 ( .A1(n725), .A2(KEYINPUT116), .ZN(n662) );
  NAND2_X1 U721 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U722 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U723 ( .A1(n667), .A2(n666), .ZN(n669) );
  XNOR2_X1 U724 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n668) );
  XNOR2_X1 U725 ( .A(n669), .B(n668), .ZN(G75) );
  NAND2_X1 U726 ( .A1(n705), .A2(G475), .ZN(n673) );
  XOR2_X1 U727 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n670) );
  XNOR2_X1 U728 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U729 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U730 ( .A1(n674), .A2(n716), .ZN(n675) );
  XNOR2_X1 U731 ( .A(n675), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U732 ( .A1(n705), .A2(G210), .ZN(n680) );
  XOR2_X1 U733 ( .A(KEYINPUT86), .B(KEYINPUT54), .Z(n677) );
  XNOR2_X1 U734 ( .A(n677), .B(KEYINPUT55), .ZN(n678) );
  XNOR2_X1 U735 ( .A(n676), .B(n678), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U737 ( .A1(n681), .A2(n716), .ZN(n683) );
  XNOR2_X1 U738 ( .A(KEYINPUT118), .B(KEYINPUT56), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n683), .B(n682), .ZN(G51) );
  XOR2_X1 U740 ( .A(G101), .B(n684), .Z(G3) );
  NAND2_X1 U741 ( .A1(n686), .A2(n696), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n685), .B(G104), .ZN(G6) );
  XOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n688) );
  NAND2_X1 U744 ( .A1(n686), .A2(n699), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U746 ( .A(G107), .B(n689), .ZN(G9) );
  XOR2_X1 U747 ( .A(G110), .B(n690), .Z(G12) );
  XOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .Z(n692) );
  NAND2_X1 U749 ( .A1(n693), .A2(n699), .ZN(n691) );
  XNOR2_X1 U750 ( .A(n692), .B(n691), .ZN(G30) );
  NAND2_X1 U751 ( .A1(n693), .A2(n696), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n694), .B(KEYINPUT110), .ZN(n695) );
  XNOR2_X1 U753 ( .A(G146), .B(n695), .ZN(G48) );
  NAND2_X1 U754 ( .A1(n698), .A2(n696), .ZN(n697) );
  XNOR2_X1 U755 ( .A(n697), .B(G113), .ZN(G15) );
  XOR2_X1 U756 ( .A(G116), .B(KEYINPUT111), .Z(n701) );
  NAND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(G18) );
  XNOR2_X1 U759 ( .A(G125), .B(n702), .ZN(n703) );
  XNOR2_X1 U760 ( .A(n703), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U761 ( .A(G134), .B(n704), .ZN(G36) );
  NAND2_X1 U762 ( .A1(n711), .A2(G469), .ZN(n709) );
  XOR2_X1 U763 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n716), .A2(n710), .ZN(G54) );
  NAND2_X1 U766 ( .A1(n711), .A2(G217), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n712), .B(KEYINPUT120), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n716), .A2(n715), .ZN(G66) );
  XOR2_X1 U769 ( .A(n717), .B(KEYINPUT122), .Z(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n720), .B(G101), .ZN(n722) );
  NOR2_X1 U772 ( .A1(n725), .A2(G898), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U774 ( .A(KEYINPUT123), .B(n723), .Z(n732) );
  NAND2_X1 U775 ( .A1(n375), .A2(n725), .ZN(n730) );
  XOR2_X1 U776 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n727) );
  NAND2_X1 U777 ( .A1(G224), .A2(G953), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U779 ( .A1(n728), .A2(G898), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(G69) );
  XNOR2_X1 U782 ( .A(n733), .B(KEYINPUT124), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n738), .B(n741), .ZN(n739) );
  XNOR2_X1 U786 ( .A(KEYINPUT125), .B(n739), .ZN(n740) );
  NOR2_X1 U787 ( .A1(G953), .A2(n740), .ZN(n745) );
  XNOR2_X1 U788 ( .A(G227), .B(n741), .ZN(n743) );
  NAND2_X1 U789 ( .A1(G900), .A2(G953), .ZN(n742) );
  NOR2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U791 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U792 ( .A(KEYINPUT126), .B(n746), .ZN(G72) );
  XNOR2_X1 U793 ( .A(G131), .B(n747), .ZN(G33) );
  XOR2_X1 U794 ( .A(G143), .B(n748), .Z(G45) );
  XNOR2_X1 U795 ( .A(n749), .B(G122), .ZN(G24) );
  XNOR2_X1 U796 ( .A(G140), .B(n750), .ZN(G42) );
  XOR2_X1 U797 ( .A(G137), .B(n751), .Z(n752) );
  XNOR2_X1 U798 ( .A(KEYINPUT127), .B(n752), .ZN(G39) );
endmodule

