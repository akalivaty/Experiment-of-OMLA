//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n208), .B(new_n211), .C1(new_n212), .C2(KEYINPUT2), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n208), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT78), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G134gat), .ZN(new_n227));
  INV_X1    g026(.A(G134gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G127gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n225), .A2(KEYINPUT1), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n240), .A3(KEYINPUT3), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n213), .A2(new_n221), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n224), .A2(new_n239), .A3(new_n241), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n230), .A2(new_n238), .A3(KEYINPUT72), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT72), .B1(new_n230), .B2(new_n238), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n242), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n230), .A2(new_n238), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n242), .A2(new_n252), .A3(KEYINPUT79), .A4(new_n247), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n213), .A2(new_n230), .A3(new_n221), .A4(new_n238), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(KEYINPUT4), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n245), .B(new_n246), .C1(new_n251), .C2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n222), .A2(new_n239), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n255), .ZN(new_n261));
  INV_X1    g060(.A(new_n246), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n239), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n230), .A2(new_n238), .A3(KEYINPUT72), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n247), .B1(new_n268), .B2(new_n222), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n242), .A2(new_n252), .A3(KEYINPUT4), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n245), .A2(new_n269), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n207), .B1(new_n264), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(new_n207), .A3(new_n272), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n273), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT81), .B1(new_n273), .B2(KEYINPUT6), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n272), .ZN(new_n283));
  INV_X1    g082(.A(new_n207), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT6), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n273), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT87), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n278), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  AND2_X1   g090(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n294), .A2(new_n299), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  AND2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  AOI211_X1 g110(.A(new_n305), .B(new_n306), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  INV_X1    g113(.A(new_n311), .ZN(new_n315));
  NOR3_X1   g114(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n316));
  OAI22_X1  g115(.A1(new_n315), .A2(new_n316), .B1(new_n308), .B2(new_n309), .ZN(new_n317));
  NOR2_X1   g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n300), .A2(new_n302), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n305), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT64), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT64), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n322), .B(new_n305), .C1(new_n317), .C2(new_n319), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n312), .A3(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n314), .A2(new_n321), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT71), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n306), .B1(new_n327), .B2(KEYINPUT26), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(KEYINPUT26), .B2(new_n327), .ZN(new_n329));
  OR2_X1    g128(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT27), .B(G183gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT28), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT70), .A4(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n339));
  AND2_X1   g138(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT68), .B1(new_n291), .B2(KEYINPUT27), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n330), .B2(new_n331), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n295), .B(new_n329), .C1(new_n338), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  INV_X1    g146(.A(G226gat), .ZN(new_n348));
  INV_X1    g147(.A(G233gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n345), .A3(new_n350), .ZN(new_n353));
  XNOR2_X1  g152(.A(G197gat), .B(G204gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT22), .ZN(new_n355));
  INV_X1    g154(.A(G211gat), .ZN(new_n356));
  INV_X1    g155(.A(G218gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G211gat), .B(G218gat), .Z(new_n360));
  OR2_X1    g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT76), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n352), .B(new_n353), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT29), .B(new_n350), .C1(new_n326), .C2(new_n345), .ZN(new_n367));
  INV_X1    g166(.A(new_n353), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G8gat), .B(G36gat), .Z(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G64gat), .ZN(new_n372));
  INV_X1    g171(.A(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n365), .B2(new_n369), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT30), .B1(new_n380), .B2(KEYINPUT77), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n369), .A3(new_n374), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n290), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n347), .B1(new_n363), .B2(new_n364), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n242), .B1(new_n386), .B2(new_n243), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n244), .A2(new_n347), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n366), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(G228gat), .B(G233gat), .C1(new_n387), .C2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n361), .A2(new_n362), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n347), .A3(new_n222), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n223), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT82), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n366), .A2(new_n388), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n399), .A3(new_n223), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(new_n392), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n392), .B1(new_n390), .B2(new_n401), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n405), .B(G22gat), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n403), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n401), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n391), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n410), .B2(new_n402), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT33), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n346), .A2(new_n268), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n326), .A2(new_n345), .A3(new_n250), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G227gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n349), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT73), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n326), .A2(new_n250), .A3(new_n345), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n250), .B1(new_n326), .B2(new_n345), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT73), .B(new_n420), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n415), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT74), .B(G15gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G43gat), .ZN(new_n428));
  XOR2_X1   g227(.A(G71gat), .B(G99gat), .Z(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n418), .A2(KEYINPUT34), .A3(new_n420), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT34), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n422), .A2(new_n423), .ZN(new_n435));
  INV_X1    g234(.A(new_n420), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n424), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n431), .A2(KEYINPUT33), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT32), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n432), .A2(new_n438), .A3(new_n444), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n433), .A2(new_n437), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n430), .B1(new_n442), .B2(new_n415), .ZN(new_n447));
  INV_X1    g246(.A(new_n443), .ZN(new_n448));
  AOI211_X1 g247(.A(new_n414), .B(new_n448), .C1(new_n441), .C2(new_n424), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n413), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n202), .B1(new_n385), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n445), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(new_n412), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n454), .A2(KEYINPUT35), .A3(new_n456), .A4(new_n384), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n447), .A2(new_n449), .A3(new_n446), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n438), .B1(new_n432), .B2(new_n444), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT75), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n408), .B2(new_n411), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n410), .A2(new_n406), .A3(new_n402), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT83), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n455), .B2(new_n383), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n453), .A2(KEYINPUT75), .A3(KEYINPUT36), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n462), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n245), .A2(new_n269), .A3(new_n270), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n262), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n260), .A2(new_n246), .A3(new_n255), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT39), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n476), .A3(new_n262), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n207), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(KEYINPUT40), .A3(new_n207), .A4(new_n477), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n480), .A2(new_n481), .A3(new_n274), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n383), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n413), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n370), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT37), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n374), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n281), .B1(new_n279), .B2(new_n280), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n288), .ZN(new_n490));
  AOI221_X4 g289(.A(new_n277), .B1(new_n488), .B2(KEYINPUT38), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT38), .B1(new_n487), .B2(KEYINPUT84), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n375), .B1(new_n370), .B2(new_n485), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n365), .A2(new_n369), .A3(new_n494), .A4(KEYINPUT37), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT86), .A4(new_n495), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n380), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n484), .B1(new_n491), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n452), .B(new_n457), .C1(new_n471), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504));
  INV_X1    g303(.A(G71gat), .ZN(new_n505));
  INV_X1    g304(.A(G78gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT97), .ZN(new_n508));
  XOR2_X1   g307(.A(G57gat), .B(G64gat), .Z(new_n509));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n504), .C1(new_n505), .C2(new_n506), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n514), .B(new_n515), .Z(new_n516));
  OR2_X1    g315(.A1(new_n516), .A2(KEYINPUT21), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n517), .B(new_n518), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT16), .A3(new_n522), .ZN(new_n523));
  OAI221_X1 g322(.A(new_n523), .B1(KEYINPUT94), .B2(G8gat), .C1(new_n522), .C2(new_n521), .ZN(new_n524));
  NAND2_X1  g323(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(KEYINPUT21), .B2(new_n516), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(new_n291), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT98), .ZN(new_n529));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(new_n356), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n530), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n529), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n533), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n520), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(new_n533), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n519), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(G29gat), .A2(G36gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT14), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT92), .Z(new_n546));
  XOR2_X1   g345(.A(KEYINPUT90), .B(G36gat), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G29gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT93), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT91), .B(G50gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(G43gat), .ZN(new_n552));
  INV_X1    g351(.A(G43gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G50gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(G50gat), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n556), .A2(new_n554), .A3(new_n550), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n548), .B2(KEYINPUT93), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n546), .A2(new_n549), .A3(new_n555), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n548), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n560), .B2(new_n545), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT17), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n559), .B2(new_n561), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT7), .ZN(new_n568));
  INV_X1    g367(.A(G99gat), .ZN(new_n569));
  INV_X1    g368(.A(G106gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT8), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n568), .B(new_n571), .C1(G85gat), .C2(G92gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT100), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n572), .B(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(new_n573), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT101), .B1(new_n566), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n562), .B2(new_n577), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT101), .ZN(new_n581));
  INV_X1    g380(.A(new_n577), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n581), .B(new_n582), .C1(new_n563), .C2(new_n565), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G190gat), .ZN(new_n585));
  INV_X1    g384(.A(G190gat), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n578), .A2(new_n586), .A3(new_n580), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n357), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(G218gat), .A3(new_n587), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n503), .A2(new_n543), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n526), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n563), .B2(new_n565), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n562), .A2(new_n526), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n604), .A2(KEYINPUT95), .A3(KEYINPUT18), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n562), .B(new_n526), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n605), .B(KEYINPUT13), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n602), .A2(new_n603), .A3(new_n605), .A4(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n606), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT89), .ZN(new_n616));
  XOR2_X1   g415(.A(G113gat), .B(G141gat), .Z(new_n617));
  XNOR2_X1  g416(.A(G169gat), .B(G197gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n615), .A2(KEYINPUT89), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n349), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n572), .B(new_n574), .Z(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n516), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n516), .B2(new_n577), .ZN(new_n633));
  INV_X1    g432(.A(new_n516), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n582), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT10), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n516), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n628), .A3(new_n635), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n309), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n638), .B2(new_n639), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n626), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n600), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n600), .A2(KEYINPUT104), .A3(new_n649), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n455), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT16), .ZN(new_n658));
  INV_X1    g457(.A(G8gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n383), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n661), .A2(new_n657), .A3(new_n662), .ZN(new_n667));
  INV_X1    g466(.A(new_n654), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n668), .B2(new_n384), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n665), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(G1325gat));
  INV_X1    g469(.A(new_n453), .ZN(new_n671));
  AOI21_X1  g470(.A(G15gat), .B1(new_n654), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n462), .A2(new_n470), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n674), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n468), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AND2_X1   g477(.A1(new_n502), .A2(new_n599), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n539), .A2(new_n542), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n626), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n681), .A3(new_n647), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n682), .A2(G29gat), .A3(new_n456), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(G29gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n471), .A2(new_n501), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n452), .A2(new_n457), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT108), .B(new_n599), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n502), .A2(KEYINPUT108), .A3(KEYINPUT44), .A4(new_n599), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n647), .B(KEYINPUT107), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n680), .A2(new_n626), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT109), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n691), .A2(new_n695), .A3(new_n698), .A4(new_n692), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n456), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n685), .B1(new_n686), .B2(new_n700), .ZN(G1328gat));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT110), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n682), .A2(new_n547), .A3(new_n384), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(KEYINPUT110), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n547), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n384), .B1(new_n697), .B2(new_n699), .ZN(new_n708));
  OAI221_X1 g507(.A(new_n706), .B1(new_n703), .B2(new_n704), .C1(new_n707), .C2(new_n708), .ZN(G1329gat));
  NOR3_X1   g508(.A1(new_n682), .A2(G43gat), .A3(new_n453), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G43gat), .B1(new_n696), .B2(new_n673), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(KEYINPUT47), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n699), .ZN(new_n714));
  INV_X1    g513(.A(new_n673), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n710), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n717), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g517(.A(new_n551), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n696), .B2(new_n413), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n551), .B(new_n468), .C1(new_n682), .C2(KEYINPUT112), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n682), .A2(KEYINPUT112), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n720), .B(KEYINPUT48), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n468), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n719), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT113), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(new_n723), .C1(new_n726), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n543), .A2(new_n599), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n626), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n503), .A3(new_n693), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n455), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  INV_X1    g536(.A(new_n735), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n383), .A2(KEYINPUT114), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n383), .A2(KEYINPUT114), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n738), .B2(new_n673), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n735), .A2(new_n505), .A3(new_n671), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n468), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g551(.A1(new_n691), .A2(new_n692), .ZN(new_n753));
  INV_X1    g552(.A(new_n626), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n680), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n648), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756), .B2(new_n456), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n679), .A2(new_n755), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT115), .Z(new_n761));
  INV_X1    g560(.A(G85gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n762), .A3(new_n648), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n763), .B2(new_n456), .ZN(G1336gat));
  INV_X1    g563(.A(new_n741), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n760), .A2(new_n373), .A3(new_n694), .A4(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n756), .B2(new_n741), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G92gat), .B1(new_n756), .B2(new_n384), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(new_n768), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n756), .B2(new_n673), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n761), .A2(new_n569), .A3(new_n648), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n453), .ZN(G1338gat));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n570), .A3(new_n412), .A4(new_n694), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G106gat), .B1(new_n756), .B2(new_n413), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND4_X1   g580(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n780), .ZN(new_n782));
  INV_X1    g581(.A(new_n468), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n756), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n781), .A2(new_n782), .B1(new_n778), .B2(new_n785), .ZN(G1339gat));
  OR3_X1    g585(.A1(new_n636), .A2(new_n637), .A3(new_n629), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(KEYINPUT54), .A3(new_n638), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n629), .C1(new_n636), .C2(new_n637), .ZN(new_n790));
  INV_X1    g589(.A(new_n643), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n788), .A2(new_n792), .A3(KEYINPUT55), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n644), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT117), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n795), .A2(new_n799), .A3(new_n644), .A4(new_n796), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n754), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n604), .A2(new_n605), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n607), .A2(new_n608), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n621), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n615), .B2(new_n622), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n648), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n599), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n599), .A2(new_n798), .A3(new_n800), .A4(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n543), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n733), .A2(new_n647), .A3(new_n626), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n813), .A2(new_n456), .A3(new_n451), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n741), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n233), .A3(new_n754), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n813), .A2(new_n468), .A3(new_n453), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n765), .A2(new_n456), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819), .B2(new_n626), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(G1340gat));
  OAI21_X1  g620(.A(G120gat), .B1(new_n819), .B2(new_n693), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n814), .A2(new_n231), .A3(new_n648), .A4(new_n741), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(KEYINPUT118), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n815), .B2(new_n680), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n819), .A2(new_n226), .A3(new_n543), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(G1342gat));
  INV_X1    g630(.A(new_n599), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n383), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n228), .A3(new_n833), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT56), .Z(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n819), .B2(new_n832), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1343gat));
  INV_X1    g636(.A(new_n797), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n754), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  OR3_X1    g639(.A1(new_n805), .A2(new_n647), .A3(KEYINPUT119), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT119), .B1(new_n805), .B2(new_n647), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n797), .A2(new_n626), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT120), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n846), .A3(new_n832), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n680), .B1(new_n847), .B2(new_n809), .ZN(new_n848));
  INV_X1    g647(.A(new_n812), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n468), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n818), .A2(new_n673), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n811), .A2(new_n812), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n412), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n851), .A2(new_n754), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT121), .B1(new_n853), .B2(new_n455), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n859), .B(new_n456), .C1(new_n811), .C2(new_n812), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n715), .A2(new_n413), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT122), .Z(new_n863));
  NAND2_X1  g662(.A1(new_n754), .A2(new_n214), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT123), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n861), .A2(new_n741), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n861), .A2(new_n863), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n765), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n216), .A3(new_n648), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n647), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n216), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n813), .B2(new_n413), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n599), .A2(new_n838), .A3(new_n806), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n680), .B1(new_n847), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n854), .B(new_n468), .C1(new_n881), .C2(new_n849), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n879), .A2(new_n648), .A3(new_n852), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n875), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n874), .B1(new_n878), .B2(new_n884), .ZN(G1345gat));
  NOR3_X1   g684(.A1(new_n876), .A2(new_n209), .A3(new_n543), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n873), .A2(new_n680), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n209), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n876), .B2(new_n832), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n833), .A2(new_n210), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n872), .B2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n384), .A2(new_n455), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n817), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n626), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n813), .A2(new_n455), .A3(new_n741), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n308), .A3(new_n454), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n626), .B2(new_n896), .ZN(G1348gat));
  OAI21_X1  g696(.A(G176gat), .B1(new_n893), .B2(new_n693), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n895), .A2(new_n309), .A3(new_n454), .A4(new_n648), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  NOR2_X1   g702(.A1(new_n813), .A2(new_n453), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(new_n680), .A3(new_n783), .A4(new_n892), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G183gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n895), .A2(new_n454), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n680), .A2(new_n333), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n906), .B(new_n911), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n893), .B2(new_n832), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n895), .A2(new_n599), .A3(new_n332), .A4(new_n454), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n914), .A2(new_n916), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(G1351gat));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n895), .A2(new_n923), .A3(new_n754), .A4(new_n862), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT127), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n673), .A2(new_n892), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n879), .A2(new_n882), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n626), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(G1352gat));
  AND2_X1   g728(.A1(new_n895), .A2(new_n862), .ZN(new_n930));
  INV_X1    g729(.A(G204gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n648), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  OAI21_X1  g732(.A(G204gat), .B1(new_n927), .B2(new_n693), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n930), .A2(new_n935), .A3(new_n931), .A4(new_n648), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n930), .A2(new_n356), .A3(new_n680), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n879), .A2(new_n680), .A3(new_n882), .A4(new_n926), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  NAND3_X1  g742(.A1(new_n930), .A2(new_n357), .A3(new_n599), .ZN(new_n944));
  OAI21_X1  g743(.A(G218gat), .B1(new_n927), .B2(new_n832), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


