//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n188), .A2(KEYINPUT68), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(KEYINPUT68), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT65), .A2(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT65), .A2(G134), .ZN(new_n192));
  AOI21_X1  g006(.A(G137), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G134), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT66), .A3(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(G131), .B1(new_n193), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G137), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n195), .A2(KEYINPUT11), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n191), .A2(new_n206), .A3(new_n192), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n211), .A2(new_n213), .B1(new_n215), .B2(G128), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT67), .A3(new_n211), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n216), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n209), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT0), .A4(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n214), .A2(G143), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n212), .A2(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n210), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n224), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n191), .A2(new_n206), .A3(new_n192), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n201), .A2(new_n203), .ZN(new_n236));
  OAI21_X1  g050(.A(G131), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n208), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n189), .B(new_n190), .C1(new_n223), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n216), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT67), .B1(new_n220), .B2(new_n211), .ZN(new_n241));
  AND4_X1   g055(.A1(KEYINPUT67), .A2(new_n211), .A3(new_n213), .A4(new_n215), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n208), .A3(new_n200), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n226), .A2(new_n227), .A3(new_n225), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n213), .A2(new_n215), .B1(KEYINPUT0), .B2(G128), .ZN(new_n246));
  INV_X1    g060(.A(new_n233), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n208), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n205), .B1(new_n204), .B2(new_n207), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n244), .A2(new_n251), .A3(KEYINPUT68), .A4(new_n188), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n239), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G119), .ZN(new_n256));
  INV_X1    g070(.A(G119), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT69), .A3(G116), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G119), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT2), .B(G113), .Z(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  INV_X1    g078(.A(new_n262), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n244), .A3(new_n251), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  INV_X1    g089(.A(new_n271), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n244), .A2(new_n251), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n262), .B1(new_n277), .B2(KEYINPUT72), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n244), .A2(new_n251), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT28), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n262), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n266), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n276), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n263), .A2(new_n273), .A3(new_n286), .A4(new_n264), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n275), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n265), .B1(new_n239), .B2(new_n252), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT31), .B1(new_n289), .B2(new_n272), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT70), .B(KEYINPUT31), .C1(new_n289), .C2(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n298), .B(new_n187), .C1(new_n288), .C2(new_n294), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G472), .ZN(new_n301));
  INV_X1    g115(.A(new_n284), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n278), .A2(new_n280), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n271), .B(new_n302), .C1(new_n303), .C2(KEYINPUT28), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n263), .A2(new_n266), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n304), .B(new_n305), .C1(new_n271), .C2(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n281), .A2(new_n284), .A3(new_n276), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n301), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n187), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n275), .A2(new_n285), .A3(new_n287), .ZN(new_n313));
  INV_X1    g127(.A(new_n294), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(KEYINPUT32), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n300), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT9), .B(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  INV_X1    g136(.A(G227), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n327));
  INV_X1    g141(.A(G107), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G104), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(G104), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(KEYINPUT82), .ZN(new_n331));
  INV_X1    g145(.A(G104), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G101), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n332), .B2(G107), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(KEYINPUT3), .A3(G104), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(KEYINPUT79), .A2(G101), .ZN(new_n341));
  NOR2_X1   g155(.A1(KEYINPUT79), .A2(G101), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND4_X1   g157(.A1(KEYINPUT80), .A2(new_n340), .A3(new_n343), .A4(new_n333), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT80), .B1(new_n345), .B2(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n327), .B1(new_n347), .B2(new_n222), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n328), .A2(KEYINPUT3), .A3(G104), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT3), .B1(new_n328), .B2(G104), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n333), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n349), .B1(new_n352), .B2(G101), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n344), .B2(new_n346), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(G101), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n248), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n358));
  INV_X1    g172(.A(new_n343), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n358), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n345), .A2(KEYINPUT80), .A3(new_n343), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(KEYINPUT10), .A3(new_n243), .A4(new_n336), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n357), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n249), .A2(new_n250), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(KEYINPUT84), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n348), .A2(new_n357), .A3(new_n363), .A4(new_n365), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n326), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n326), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n375));
  NAND2_X1  g189(.A1(new_n347), .A2(new_n222), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n243), .A3(new_n336), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n365), .B(new_n381), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n374), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n320), .B(new_n321), .C1(new_n373), .C2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n320), .A2(new_n321), .ZN(new_n386));
  INV_X1    g200(.A(new_n374), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n372), .B1(new_n379), .B2(new_n382), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n371), .A2(new_n387), .B1(new_n325), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n386), .B1(new_n389), .B2(G469), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G214), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G210), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n354), .A2(new_n262), .A3(new_n356), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n260), .A2(new_n261), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT5), .A4(new_n259), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n255), .A2(KEYINPUT5), .A3(G119), .ZN(new_n399));
  INV_X1    g213(.A(G113), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n362), .A2(new_n397), .A3(new_n336), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G122), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT6), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n396), .A2(new_n403), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n404), .B(KEYINPUT85), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n411));
  INV_X1    g225(.A(G224), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n234), .A2(new_n414), .A3(G125), .ZN(new_n415));
  INV_X1    g229(.A(G125), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n416), .B(new_n240), .C1(new_n241), .C2(new_n242), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n234), .B2(G125), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n418), .A2(new_n413), .A3(new_n419), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n410), .A2(new_n411), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n404), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n397), .A2(new_n402), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n347), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n403), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  OAI22_X1  g243(.A1(new_n418), .A2(new_n419), .B1(new_n429), .B2(new_n413), .ZN(new_n430));
  INV_X1    g244(.A(new_n419), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n413), .A2(new_n429), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n417), .A3(new_n415), .A4(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n428), .A2(new_n405), .A3(new_n430), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n321), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n395), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n421), .A2(new_n420), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n405), .A2(KEYINPUT6), .B1(new_n407), .B2(new_n408), .ZN(new_n438));
  INV_X1    g252(.A(new_n411), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n433), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(new_n427), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n442), .B2(new_n405), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n443), .A3(new_n394), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n393), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n446));
  XOR2_X1   g260(.A(G116), .B(G122), .Z(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  XNOR2_X1  g262(.A(G116), .B(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n328), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n212), .A2(G128), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n210), .A2(G143), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n452), .A2(new_n453), .ZN(new_n457));
  OAI21_X1  g271(.A(G134), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n191), .A2(new_n192), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n452), .A2(new_n455), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n451), .A2(new_n458), .A3(KEYINPUT90), .A4(new_n461), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n459), .B(new_n460), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n255), .A2(KEYINPUT14), .A3(G122), .ZN(new_n467));
  OAI211_X1 g281(.A(G107), .B(new_n467), .C1(new_n447), .C2(KEYINPUT14), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n450), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G217), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n318), .A2(new_n471), .A3(G953), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n464), .A2(new_n465), .A3(new_n469), .A4(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n446), .B1(new_n476), .B2(new_n321), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT91), .B(G902), .C1(new_n474), .C2(new_n475), .ZN(new_n478));
  INV_X1    g292(.A(G478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT15), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G237), .ZN(new_n483));
  INV_X1    g297(.A(G953), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(G214), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n212), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT18), .A2(G131), .ZN(new_n489));
  XNOR2_X1  g303(.A(G125), .B(G140), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n490), .A2(new_n214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n214), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n488), .A2(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n487), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT18), .A3(G131), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n332), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n205), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n490), .A2(KEYINPUT16), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n416), .A2(KEYINPUT16), .A3(G140), .ZN(new_n505));
  AOI21_X1  g319(.A(G146), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(G146), .A3(new_n505), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n494), .A2(KEYINPUT17), .A3(G131), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n496), .B(new_n498), .C1(new_n503), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n502), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n498), .B1(new_n513), .B2(new_n496), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n321), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G475), .ZN(new_n516));
  INV_X1    g330(.A(new_n508), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n501), .B2(new_n499), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n490), .B2(KEYINPUT89), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT19), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT19), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n490), .B2(new_n519), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n521), .B(new_n214), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n518), .A2(new_n524), .B1(new_n495), .B2(new_n493), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n511), .B1(new_n525), .B2(new_n498), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  NOR2_X1   g341(.A1(G475), .A2(G902), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(G234), .A2(G237), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n532), .A2(G952), .A3(new_n484), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(G902), .A3(G953), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT92), .Z(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n476), .A2(new_n321), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n480), .ZN(new_n539));
  NOR4_X1   g353(.A1(new_n482), .A2(new_n531), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n319), .A2(new_n391), .A3(new_n445), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(G217), .A2(G902), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n471), .B2(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT74), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n257), .A2(G128), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n257), .A2(G128), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT24), .B(G110), .Z(new_n549));
  NAND3_X1  g363(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(new_n547), .C1(new_n545), .C2(KEYINPUT23), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n548), .A2(new_n549), .B1(G110), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n508), .A3(new_n492), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(G110), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT75), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n549), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n517), .B2(new_n506), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n484), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n553), .B(new_n562), .C1(new_n555), .C2(new_n557), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n321), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n544), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n564), .A2(new_n565), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n544), .A2(G902), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT78), .Z(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n317), .A2(new_n541), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(new_n359), .ZN(G3));
  OAI21_X1  g394(.A(new_n321), .B1(new_n288), .B2(new_n294), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n296), .A2(new_n582), .A3(new_n299), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n364), .A2(KEYINPUT84), .A3(new_n366), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT84), .B1(new_n364), .B2(new_n366), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n372), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n384), .B1(new_n586), .B2(new_n325), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n587), .A2(G469), .A3(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n371), .A2(new_n387), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n388), .A2(new_n325), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(G469), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n386), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n319), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NOR4_X1   g408(.A1(new_n583), .A2(new_n594), .A3(new_n577), .A4(new_n537), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n444), .A2(KEYINPUT93), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n393), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n436), .A2(KEYINPUT93), .A3(new_n444), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n538), .A2(KEYINPUT91), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n476), .A2(new_n446), .A3(new_n321), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n479), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n476), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n479), .A2(G902), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT33), .B(new_n475), .C1(new_n474), .C2(KEYINPUT95), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n474), .A2(KEYINPUT95), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n526), .A2(new_n528), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT20), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n602), .A2(new_n608), .B1(new_n612), .B2(new_n516), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n599), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n595), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n539), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n600), .A2(new_n480), .A3(new_n601), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n531), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n599), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n595), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  AND3_X1   g440(.A1(new_n296), .A2(new_n582), .A3(new_n299), .ZN(new_n627));
  INV_X1    g441(.A(new_n594), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n558), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n575), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n572), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n610), .A2(new_n611), .B1(G475), .B2(new_n515), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n619), .A3(new_n620), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n633), .A2(new_n635), .A3(new_n537), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n627), .A2(new_n628), .A3(new_n445), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n533), .B1(new_n535), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AND4_X1   g456(.A1(new_n598), .A2(new_n597), .A3(new_n621), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n317), .A2(new_n643), .A3(new_n628), .A4(new_n632), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n594), .B1(new_n300), .B2(new_n316), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n647), .A2(KEYINPUT96), .A3(new_n632), .A4(new_n643), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XOR2_X1   g464(.A(new_n641), .B(KEYINPUT39), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n628), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n306), .A2(new_n271), .ZN(new_n655));
  INV_X1    g469(.A(new_n283), .ZN(new_n656));
  INV_X1    g470(.A(new_n266), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n658), .B2(new_n276), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n301), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n315), .B2(KEYINPUT32), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n300), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n436), .A2(new_n444), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n531), .B1(new_n482), .B2(new_n539), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n665), .A2(new_n393), .A3(new_n632), .A4(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n653), .A2(new_n654), .A3(new_n662), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  NAND2_X1  g483(.A1(new_n602), .A2(new_n608), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n670), .A2(new_n531), .A3(new_n642), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n598), .A3(new_n597), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(KEYINPUT98), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n647), .A2(new_n673), .A3(new_n632), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  OAI21_X1  g490(.A(G469), .B1(new_n587), .B2(G902), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n385), .A3(KEYINPUT99), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n679), .B(G469), .C1(new_n587), .C2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n319), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n537), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n577), .B1(new_n300), .B2(new_n316), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n615), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n684), .A3(new_n623), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND4_X1  g503(.A1(new_n681), .A2(new_n319), .A3(new_n598), .A4(new_n597), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n317), .A3(new_n636), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n599), .A2(new_n694), .A3(new_n666), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n694), .B1(new_n599), .B2(new_n666), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n312), .B1(new_n313), .B2(new_n290), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n582), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n581), .A2(KEYINPUT100), .A3(G472), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n683), .A3(new_n578), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT102), .B(G122), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G24));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n701), .ZN(new_n706));
  INV_X1    g520(.A(new_n698), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n632), .A3(new_n671), .A4(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n690), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n416), .ZN(G27));
  AND2_X1   g524(.A1(new_n436), .A2(new_n444), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n392), .A3(new_n613), .A4(new_n642), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n594), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n295), .A2(new_n297), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n577), .B1(new_n316), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n594), .A2(new_n712), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n317), .A2(new_n719), .A3(KEYINPUT103), .A4(new_n578), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n684), .B2(new_n719), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT104), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n317), .A2(new_n719), .A3(new_n578), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n713), .A4(new_n720), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n718), .B1(new_n723), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n205), .ZN(G33));
  AND3_X1   g544(.A1(new_n436), .A2(new_n392), .A3(new_n444), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n732), .A2(new_n622), .A3(new_n577), .A4(new_n641), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n647), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  NAND2_X1  g549(.A1(new_n670), .A2(new_n634), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(KEYINPUT43), .Z(new_n737));
  AND3_X1   g551(.A1(new_n583), .A2(KEYINPUT105), .A3(new_n632), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT105), .B1(new_n583), .B2(new_n632), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n389), .A2(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n389), .A2(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(G469), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT46), .B1(new_n745), .B2(new_n592), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n588), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n592), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n749), .A2(new_n319), .A3(new_n651), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n740), .A2(new_n741), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n742), .A2(new_n750), .A3(new_n731), .A4(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT106), .B(G137), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G39));
  NOR3_X1   g568(.A1(new_n317), .A2(new_n578), .A3(new_n712), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n749), .A2(new_n319), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n319), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  INV_X1    g577(.A(new_n681), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT49), .ZN(new_n765));
  INV_X1    g579(.A(new_n665), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n578), .A2(new_n319), .A3(new_n392), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n766), .A2(new_n736), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n662), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n764), .A2(KEYINPUT49), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n765), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n533), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n682), .A2(new_n772), .A3(new_n732), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n578), .A3(new_n769), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n634), .A3(new_n602), .A4(new_n608), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n773), .A2(new_n737), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n633), .B(new_n698), .C1(new_n700), .C2(new_n701), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n702), .A2(new_n578), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n737), .A2(new_n533), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n682), .A2(new_n766), .A3(new_n392), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n758), .B(new_n760), .C1(new_n319), .C2(new_n764), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n782), .A2(new_n783), .A3(new_n732), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n792), .A3(KEYINPUT51), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n784), .A2(new_n691), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(G952), .A3(new_n484), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n777), .A2(new_n716), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT48), .Z(new_n798));
  AOI211_X1 g612(.A(new_n796), .B(new_n798), .C1(new_n613), .C2(new_n775), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n792), .A2(new_n779), .A3(new_n776), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n794), .B(new_n799), .C1(KEYINPUT51), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n723), .A2(new_n728), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n717), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n703), .A2(new_n685), .A3(new_n688), .A4(new_n692), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n482), .A2(new_n531), .A3(new_n539), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n731), .A2(new_n807), .A3(KEYINPUT107), .A4(new_n642), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT107), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n436), .A2(new_n444), .A3(new_n392), .A4(new_n642), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n635), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n317), .A3(new_n628), .A4(new_n632), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n702), .A2(new_n632), .A3(new_n719), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n734), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n577), .A2(new_n537), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n621), .A2(new_n613), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n663), .A2(new_n392), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n627), .A2(new_n628), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n579), .A2(new_n820), .A3(new_n637), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n804), .A2(new_n806), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n709), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n594), .A2(new_n632), .A3(new_n641), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n697), .A2(new_n662), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n649), .A2(new_n824), .A3(new_n675), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n709), .B1(new_n646), .B2(new_n648), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n675), .A4(new_n826), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n802), .B1(new_n823), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n579), .A2(new_n637), .A3(new_n820), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT108), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n778), .A2(new_n719), .B1(new_n647), .B2(new_n733), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n813), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT108), .B1(new_n815), .B2(new_n821), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n829), .A2(new_n830), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n729), .A2(new_n805), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n831), .A3(new_n828), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT109), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n833), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n833), .A2(new_n843), .A3(new_n845), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT109), .ZN(new_n848));
  INV_X1    g662(.A(new_n832), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n802), .B1(new_n829), .B2(new_n830), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n842), .A3(new_n822), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n845), .B1(new_n851), .B2(new_n833), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n846), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT110), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n846), .C1(new_n848), .C2(new_n852), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n801), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(G952), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n484), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT113), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n771), .B1(new_n857), .B2(new_n860), .ZN(G75));
  NAND2_X1  g675(.A1(new_n858), .A2(G953), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT115), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n321), .B1(new_n833), .B2(new_n843), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n864), .B2(G210), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n438), .A2(new_n439), .A3(new_n437), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n422), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n863), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n868), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(KEYINPUT114), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(KEYINPUT114), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G51));
  INV_X1    g687(.A(new_n863), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n833), .A2(new_n843), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n847), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n386), .B(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n587), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(KEYINPUT116), .A3(new_n878), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n745), .B(KEYINPUT117), .Z(new_n885));
  NAND2_X1  g699(.A1(new_n864), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n874), .B1(new_n884), .B2(new_n886), .ZN(G54));
  INV_X1    g701(.A(new_n526), .ZN(new_n888));
  AND2_X1   g702(.A1(KEYINPUT58), .A2(G475), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n864), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n864), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n863), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(G60));
  OR2_X1    g708(.A1(new_n606), .A2(new_n607), .ZN(new_n895));
  XNOR2_X1  g709(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n877), .A2(new_n895), .A3(new_n604), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n863), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n854), .A2(new_n856), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n604), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G63));
  XNOR2_X1  g717(.A(new_n542), .B(KEYINPUT121), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n875), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n863), .B1(new_n906), .B2(new_n573), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n630), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n906), .A2(KEYINPUT122), .A3(new_n630), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n913));
  INV_X1    g727(.A(new_n911), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n906), .B2(new_n630), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT123), .B1(new_n906), .B2(new_n573), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n875), .A2(new_n905), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n919));
  INV_X1    g733(.A(new_n573), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n917), .A2(KEYINPUT61), .A3(new_n863), .A4(new_n921), .ZN(new_n922));
  OAI22_X1  g736(.A1(new_n912), .A2(new_n913), .B1(new_n916), .B2(new_n922), .ZN(G66));
  NOR2_X1   g737(.A1(new_n805), .A2(new_n821), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(G953), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT124), .ZN(new_n926));
  OAI21_X1  g740(.A(G953), .B1(new_n536), .B2(new_n412), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n410), .B(new_n411), .C1(G898), .C2(new_n484), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G69));
  AND2_X1   g744(.A1(new_n829), .A2(new_n675), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n668), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT125), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n762), .A2(new_n752), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n652), .A2(new_n732), .A3(new_n817), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n684), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(KEYINPUT62), .B2(new_n932), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n520), .A2(new_n523), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(KEYINPUT19), .B2(new_n520), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n253), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n697), .A2(new_n716), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n750), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n931), .A2(new_n734), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n935), .A2(new_n948), .A3(new_n804), .ZN(new_n949));
  AOI21_X1  g763(.A(G953), .B1(new_n949), .B2(new_n943), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n943), .A2(G227), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n640), .B(new_n484), .C1(new_n944), .C2(new_n323), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n945), .A2(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G72));
  NAND2_X1  g767(.A1(new_n307), .A2(new_n276), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n655), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n851), .B2(new_n833), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n934), .A2(new_n939), .A3(new_n924), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n655), .B1(new_n959), .B2(new_n956), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n935), .A2(new_n948), .A3(new_n804), .A4(new_n924), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n956), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n954), .B(KEYINPUT126), .Z(new_n963));
  AOI21_X1  g777(.A(new_n874), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT127), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT127), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n958), .B(new_n960), .C1(new_n965), .C2(new_n966), .ZN(G57));
endmodule


