//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OR3_X1    g002(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT93), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NOR3_X1   g005(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT93), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n206), .A2(new_n208), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n210), .A2(KEYINPUT15), .B1(new_n203), .B2(new_n207), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n212), .A2(KEYINPUT17), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G1gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G1gat), .B2(new_n220), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(G8gat), .Z(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n211), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(new_n217), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n218), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n223), .B(G8gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT94), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n229), .B(KEYINPUT13), .Z(new_n238));
  INV_X1    g037(.A(new_n232), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n230), .A2(new_n231), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n235), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n237), .A2(new_n248), .A3(new_n241), .A4(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT64), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT24), .ZN(new_n259));
  NOR2_X1   g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(KEYINPUT23), .ZN(new_n261));
  INV_X1    g060(.A(G183gat), .ZN(new_n262));
  INV_X1    g061(.A(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT24), .A3(new_n257), .ZN(new_n265));
  INV_X1    g064(.A(new_n260), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n261), .A2(new_n265), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n269), .B(KEYINPUT65), .Z(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n266), .B2(new_n267), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n265), .A3(new_n261), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT66), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n279), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n260), .A2(KEYINPUT66), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n258), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G183gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n286), .A3(new_n263), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT28), .A3(new_n263), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n283), .A2(new_n292), .A3(KEYINPUT67), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT67), .B1(new_n283), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n276), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT1), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n297), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n300), .B(new_n276), .C1(new_n293), .C2(new_n294), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n256), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n304), .A2(KEYINPUT33), .ZN(new_n307));
  XNOR2_X1  g106(.A(G15gat), .B(G43gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G71gat), .B(G99gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n306), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n303), .A3(new_n256), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT34), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n303), .ZN(new_n318));
  AOI221_X4 g117(.A(new_n317), .B1(KEYINPUT33), .B2(new_n312), .C1(new_n318), .C2(new_n255), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n304), .B2(KEYINPUT33), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n304), .A2(new_n317), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n315), .B1(new_n324), .B2(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT31), .B(G50gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(G228gat), .ZN(new_n331));
  INV_X1    g130(.A(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G162gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT77), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT76), .B(G162gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(KEYINPUT2), .C1(new_n344), .C2(new_n335), .ZN(new_n345));
  XOR2_X1   g144(.A(G155gat), .B(G162gat), .Z(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n346), .B(new_n350), .C1(KEYINPUT2), .C2(new_n347), .ZN(new_n351));
  AND2_X1   g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT2), .ZN(new_n354));
  XNOR2_X1  g153(.A(G155gat), .B(G162gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G211gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT71), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G211gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT22), .B1(new_n365), .B2(G218gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G197gat), .B(G204gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n360), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G218gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n362), .B2(new_n364), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n367), .B(new_n359), .C1(new_n371), .C2(KEYINPUT22), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n358), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n349), .A2(new_n357), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n334), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT80), .B(new_n334), .C1(new_n375), .C2(new_n380), .ZN(new_n384));
  INV_X1    g183(.A(new_n372), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT22), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT71), .B(G211gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(new_n370), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n359), .B1(new_n388), .B2(new_n367), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n379), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n377), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT81), .B1(new_n391), .B2(new_n358), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT81), .B(new_n358), .C1(new_n373), .C2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n333), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n379), .ZN(new_n396));
  INV_X1    g195(.A(new_n376), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT82), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399));
  AOI211_X1 g198(.A(new_n399), .B(new_n376), .C1(new_n378), .C2(new_n379), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT83), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n380), .B(KEYINPUT82), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n374), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n334), .B1(new_n406), .B2(new_n393), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  AOI221_X4 g207(.A(new_n330), .B1(new_n383), .B2(new_n384), .C1(new_n402), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n330), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n402), .A2(new_n408), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n384), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n409), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n395), .A2(new_n401), .A3(KEYINPUT83), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n404), .B1(new_n403), .B2(new_n407), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n330), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n411), .A2(new_n410), .A3(new_n412), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n327), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT92), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n415), .B1(new_n409), .B2(new_n413), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n414), .A3(new_n421), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n327), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(KEYINPUT35), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT70), .B1(new_n321), .B2(new_n325), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT70), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n324), .A2(new_n319), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n316), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n431), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n327), .A2(KEYINPUT36), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n427), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT72), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n272), .A2(new_n275), .B1(new_n292), .B2(new_n283), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n283), .A2(new_n292), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n283), .A2(new_n292), .A3(KEYINPUT67), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n451), .A2(new_n452), .B1(new_n272), .B2(new_n275), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n448), .B(new_n376), .C1(new_n453), .C2(new_n446), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n447), .A2(new_n445), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n445), .A2(KEYINPUT29), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n397), .B(new_n455), .C1(new_n453), .C2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n443), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n458), .A3(new_n443), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n461), .B2(KEYINPUT30), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT73), .Z(new_n463));
  NAND2_X1  g262(.A1(new_n358), .A2(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n301), .A3(new_n378), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n300), .A2(new_n349), .A3(new_n357), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n349), .A2(new_n357), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT4), .A3(new_n300), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n472), .B(KEYINPUT78), .Z(new_n473));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n301), .A2(new_n358), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  OAI22_X1  g276(.A1(new_n471), .A2(new_n473), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n470), .A2(new_n468), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT5), .A3(new_n475), .A4(new_n465), .ZN(new_n480));
  XOR2_X1   g279(.A(G1gat), .B(G29gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G57gat), .B(G85gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND4_X1  g284(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT6), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n485), .A3(new_n480), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n478), .B2(new_n480), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT74), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n460), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n463), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n486), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n491), .B2(KEYINPUT89), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n495), .A2(new_n462), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n432), .A2(new_n435), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n504), .A2(new_n427), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n440), .A2(new_n497), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n427), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n436), .B2(new_n437), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n295), .A2(new_n456), .B1(new_n445), .B2(new_n447), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(new_n376), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n448), .B(new_n397), .C1(new_n453), .C2(new_n446), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n443), .A2(new_n513), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n517), .B(KEYINPUT88), .C1(new_n459), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n493), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n459), .A2(new_n518), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT88), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n501), .A2(new_n524), .A3(KEYINPUT90), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT90), .B1(new_n501), .B2(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n454), .A2(new_n458), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT37), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n511), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n475), .B1(new_n479), .B2(new_n465), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT39), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n485), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT40), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n476), .A2(new_n475), .A3(new_n466), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT39), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n487), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n535), .A2(KEYINPUT85), .A3(new_n539), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT85), .B1(new_n535), .B2(new_n539), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n544), .A2(new_n536), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  INV_X1    g346(.A(new_n503), .ZN(new_n548));
  NOR4_X1   g347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n510), .B1(new_n530), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n253), .B1(new_n508), .B2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G71gat), .B(G78gat), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554));
  INV_X1    g353(.A(G71gat), .ZN(new_n555));
  INV_X1    g354(.A(G78gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G57gat), .B(G64gat), .Z(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n557), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G127gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n224), .B1(new_n563), .B2(new_n562), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(new_n335), .ZN(new_n571));
  XOR2_X1   g370(.A(G183gat), .B(G211gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n574), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(G85gat), .A3(G92gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n580), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G99gat), .ZN(new_n590));
  INV_X1    g389(.A(G106gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n584), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n584), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n583), .A2(new_n587), .A3(new_n594), .A4(new_n588), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT95), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n230), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n219), .A2(new_n227), .A3(new_n596), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n579), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n600), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n601), .A2(new_n602), .A3(new_n579), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n601), .A2(new_n602), .A3(new_n579), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n607), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n577), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n596), .A2(new_n562), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n593), .A2(new_n561), .A3(new_n559), .A4(new_n595), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n619), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n620), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n617), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT97), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n491), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n491), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n551), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g441(.A(KEYINPUT16), .B(G8gat), .Z(new_n643));
  NAND4_X1  g442(.A1(new_n551), .A2(new_n503), .A3(new_n635), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n551), .A2(new_n503), .A3(new_n635), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G8gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n644), .ZN(new_n647));
  MUX2_X1   g446(.A(new_n644), .B(new_n647), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g447(.A1(new_n551), .A2(new_n635), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n436), .A2(new_n437), .ZN(new_n650));
  OAI21_X1  g449(.A(G15gat), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n432), .A2(new_n435), .A3(G15gat), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n649), .B2(new_n652), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n649), .A2(new_n427), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT43), .B(G22gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  AOI21_X1  g455(.A(new_n613), .B1(new_n508), .B2(new_n550), .ZN(new_n657));
  INV_X1    g456(.A(new_n577), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n658), .A2(new_n253), .A3(new_n632), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n213), .A3(new_n640), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n507), .A2(new_n498), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n428), .B1(new_n427), .B2(new_n327), .ZN(new_n664));
  AOI211_X1 g463(.A(KEYINPUT92), .B(new_n326), .C1(new_n425), .C2(new_n426), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n438), .B1(new_n666), .B2(KEYINPUT35), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n550), .B(new_n663), .C1(new_n667), .C2(new_n496), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n614), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(KEYINPUT44), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n670), .B(new_n659), .C1(new_n657), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n614), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n677), .A2(new_n678), .A3(new_n659), .A4(new_n670), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n675), .A2(new_n640), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n662), .B1(new_n213), .B2(new_n680), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n660), .A2(new_n214), .A3(new_n503), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  AND3_X1   g482(.A1(new_n675), .A2(new_n503), .A3(new_n679), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n214), .B2(new_n684), .ZN(G1329gat));
  OAI21_X1  g484(.A(G43gat), .B1(new_n674), .B2(new_n650), .ZN(new_n686));
  INV_X1    g485(.A(G43gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n660), .A2(new_n687), .A3(new_n505), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(KEYINPUT47), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n688), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n436), .A3(new_n437), .A4(new_n679), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(G43gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n689), .B1(new_n692), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g492(.A1(new_n427), .A2(G50gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n660), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  OAI21_X1  g495(.A(G50gat), .B1(new_n674), .B2(new_n427), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n660), .A2(new_n698), .A3(new_n694), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT48), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n675), .A2(new_n509), .A3(new_n679), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(G50gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(KEYINPUT48), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n706), .B(new_n700), .C1(new_n703), .C2(KEYINPUT48), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1331gat));
  NAND3_X1  g507(.A1(new_n615), .A2(new_n253), .A3(new_n632), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n508), .B2(new_n550), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n640), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g511(.A(new_n710), .B(KEYINPUT103), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n548), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  AND2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n714), .B2(new_n715), .ZN(G1333gat));
  OAI21_X1  g517(.A(G71gat), .B1(new_n713), .B2(new_n650), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n710), .A2(new_n505), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT104), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(G71gat), .B2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g522(.A1(new_n713), .A2(new_n427), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(new_n556), .ZN(G1335gat));
  NOR2_X1   g524(.A1(new_n658), .A2(new_n252), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n633), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n677), .A2(new_n670), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729), .B2(new_n639), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n657), .A2(new_n726), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT51), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n640), .A2(new_n585), .A3(new_n632), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n729), .B2(new_n548), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n503), .A2(new_n586), .A3(new_n632), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n735), .B(new_n736), .C1(new_n732), .C2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n731), .A2(new_n740), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n737), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n739), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n738), .B1(new_n746), .B2(new_n736), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n729), .B2(new_n650), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n505), .A2(new_n590), .A3(new_n632), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n732), .B2(new_n749), .ZN(G1338gat));
  NOR3_X1   g549(.A1(new_n427), .A2(G106gat), .A3(new_n633), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n741), .B2(new_n742), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n677), .A2(new_n509), .A3(new_n670), .A4(new_n728), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n755), .A2(KEYINPUT107), .A3(KEYINPUT53), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n755), .B2(KEYINPUT53), .ZN(new_n757));
  INV_X1    g556(.A(new_n754), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  INV_X1    g558(.A(new_n751), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n732), .B2(new_n760), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n761), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n635), .A2(new_n253), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n621), .A2(new_n622), .A3(new_n617), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT108), .ZN(new_n765));
  INV_X1    g564(.A(new_n623), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n621), .A2(new_n622), .A3(new_n767), .A4(new_n617), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT54), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n629), .B1(new_n623), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT109), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  AOI211_X1 g574(.A(new_n775), .B(KEYINPUT55), .C1(new_n769), .C2(new_n771), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n769), .A2(KEYINPUT55), .A3(new_n771), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n631), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n239), .A2(new_n240), .A3(new_n238), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n229), .B1(new_n228), .B2(new_n232), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n247), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND4_X1   g582(.A1(new_n251), .A2(new_n610), .A3(new_n612), .A4(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n777), .A2(new_n778), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n784), .B(new_n780), .C1(new_n774), .C2(new_n776), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n780), .B(new_n252), .C1(new_n774), .C2(new_n776), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n632), .A2(new_n251), .A3(new_n783), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n614), .B1(new_n791), .B2(KEYINPUT111), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n788), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n577), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g596(.A(KEYINPUT112), .B(new_n788), .C1(new_n794), .C2(new_n792), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n763), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n640), .ZN(new_n800));
  NOR4_X1   g599(.A1(new_n800), .A2(new_n503), .A3(new_n664), .A4(new_n665), .ZN(new_n801));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n252), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n639), .A2(new_n503), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n799), .A2(new_n804), .A3(new_n427), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n799), .B2(new_n427), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n505), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT114), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n252), .A2(G113gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n802), .B1(new_n809), .B2(new_n810), .ZN(G1340gat));
  AOI21_X1  g610(.A(G120gat), .B1(new_n801), .B2(new_n632), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n632), .A2(G120gat), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n809), .B2(new_n813), .ZN(G1341gat));
  OAI21_X1  g613(.A(G127gat), .B1(new_n808), .B2(new_n577), .ZN(new_n815));
  INV_X1    g614(.A(G127gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n816), .A3(new_n658), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1342gat));
  OAI21_X1  g617(.A(G134gat), .B1(new_n808), .B2(new_n613), .ZN(new_n819));
  INV_X1    g618(.A(G134gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n801), .A2(new_n820), .A3(new_n614), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT56), .Z(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(G1343gat));
  AND2_X1   g622(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n824), .A2(new_n825), .A3(new_n503), .A4(new_n439), .ZN(new_n826));
  INV_X1    g625(.A(G141gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n252), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n803), .A2(new_n650), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n799), .A2(new_n509), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n772), .A2(new_n773), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT115), .Z(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n252), .A3(new_n780), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n614), .B1(new_n835), .B2(new_n790), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n577), .B1(new_n836), .B2(new_n788), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n763), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n427), .A2(new_n831), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n829), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n253), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(G148gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n847), .A3(new_n632), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849));
  INV_X1    g648(.A(new_n786), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n577), .B1(new_n836), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n763), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n852), .B2(new_n509), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n799), .B2(new_n839), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n633), .A3(new_n829), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n847), .B1(new_n855), .B2(KEYINPUT118), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n849), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g657(.A(KEYINPUT59), .B(new_n847), .C1(new_n841), .C2(new_n632), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G1345gat));
  NAND3_X1  g659(.A1(new_n826), .A2(new_n335), .A3(new_n658), .ZN(new_n861));
  OAI21_X1  g660(.A(G155gat), .B1(new_n842), .B2(new_n577), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1346gat));
  NAND3_X1  g664(.A1(new_n826), .A2(new_n344), .A3(new_n614), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n614), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(KEYINPUT120), .ZN(new_n868));
  INV_X1    g667(.A(new_n344), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n867), .B2(KEYINPUT120), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT121), .B(new_n866), .C1(new_n868), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n640), .A2(new_n548), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n799), .A2(new_n666), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n252), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n505), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT122), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n805), .B2(new_n806), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT123), .B(new_n880), .C1(new_n805), .C2(new_n806), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n253), .A2(new_n277), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(G1348gat));
  NAND3_X1  g686(.A1(new_n877), .A2(new_n278), .A3(new_n632), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n885), .A2(new_n632), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n278), .ZN(G1349gat));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n658), .A3(new_n884), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G183gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n290), .A3(new_n658), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n895));
  NAND2_X1  g694(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n614), .A3(new_n884), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G190gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT125), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(new_n902), .A3(G190gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(KEYINPUT61), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n899), .B2(G190gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n613), .A2(G190gat), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n905), .A2(new_n906), .B1(new_n877), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n904), .A2(new_n908), .ZN(G1351gat));
  NAND2_X1  g708(.A1(new_n876), .A2(new_n650), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n830), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n252), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n854), .A2(new_n910), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n252), .A2(G197gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  INV_X1    g714(.A(G204gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n916), .A3(new_n632), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n913), .B2(new_n632), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(G1353gat));
  NAND2_X1  g719(.A1(new_n913), .A2(new_n658), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G211gat), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n911), .A2(new_n387), .A3(new_n658), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT126), .Z(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(G1354gat));
  AOI21_X1  g726(.A(G218gat), .B1(new_n911), .B2(new_n614), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n614), .A2(G218gat), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT127), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n913), .B2(new_n930), .ZN(G1355gat));
endmodule


