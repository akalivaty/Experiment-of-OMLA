//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(new_n466), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n463), .A3(G2104), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n475), .A2(G137), .A3(new_n462), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND3_X1  g055(.A1(new_n475), .A2(G2105), .A3(new_n477), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  AND2_X1   g057(.A1(G112), .A2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(G100), .B2(new_n462), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n465), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n475), .A2(new_n462), .A3(new_n477), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(G136), .B2(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n474), .A2(new_n477), .A3(new_n466), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n474), .A2(new_n477), .A3(G126), .A4(new_n466), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n462), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n492), .A2(new_n495), .A3(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .A3(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n501), .B1(new_n509), .B2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n508), .B1(new_n514), .B2(new_n503), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n504), .A2(new_n506), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n517), .B1(new_n513), .B2(new_n516), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n515), .B1(G88), .B2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n513), .A2(new_n516), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G89), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n507), .A2(new_n526), .ZN(new_n527));
  AOI211_X1 g102(.A(KEYINPUT74), .B(new_n501), .C1(new_n504), .C2(new_n506), .ZN(new_n528));
  OAI21_X1  g103(.A(G51), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n510), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n525), .A2(new_n529), .A3(new_n534), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AND3_X1   g113(.A1(new_n531), .A2(G64), .A3(new_n532), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(G651), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n523), .A2(new_n524), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n527), .A2(new_n528), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n543), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n544), .A2(new_n550), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n532), .ZN(new_n553));
  AOI21_X1  g128(.A(KEYINPUT73), .B1(new_n510), .B2(new_n512), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G56), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n503), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT75), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(new_n516), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n507), .A2(new_n570), .A3(G53), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n523), .A2(G91), .A3(new_n524), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n510), .A2(new_n512), .ZN(new_n574));
  XOR2_X1   g149(.A(KEYINPUT76), .B(G65), .Z(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n573), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G166), .ZN(G303));
  NAND2_X1  g156(.A1(new_n520), .A2(G87), .ZN(new_n582));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n553), .B2(new_n554), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G49), .B2(new_n507), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT77), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT78), .B1(new_n544), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n523), .A2(new_n593), .A3(G86), .A4(new_n524), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n574), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G48), .B2(new_n507), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n555), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n503), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n523), .A2(G85), .A3(new_n524), .ZN(new_n602));
  OAI21_X1  g177(.A(G47), .B1(new_n527), .B2(new_n528), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT79), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT79), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(G290));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n544), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n567), .A2(KEYINPUT74), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n507), .A2(new_n526), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n574), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n615), .A2(G54), .B1(G651), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n620), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g196(.A(new_n620), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g197(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g198(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g199(.A(new_n620), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NOR2_X1   g202(.A1(new_n620), .A2(G559), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n559), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT11), .Z(G282));
  INV_X1    g208(.A(new_n632), .ZN(G323));
  AND2_X1   g209(.A1(new_n487), .A2(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(KEYINPUT81), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G111), .B2(new_n462), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(KEYINPUT81), .B2(new_n636), .ZN(new_n639));
  INV_X1    g214(.A(new_n481), .ZN(new_n640));
  AOI211_X1 g215(.A(new_n635), .B(new_n639), .C1(G123), .C2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT13), .B(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n644), .A3(new_n649), .ZN(G156));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT82), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  INV_X1    g236(.A(new_n658), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT15), .B(G2435), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2438), .ZN(new_n666));
  INV_X1    g241(.A(G2427), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(G2430), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(G2430), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n651), .B1(new_n664), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n659), .A3(new_n663), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XNOR2_X1  g252(.A(G2084), .B(G2090), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  NOR2_X1   g254(.A1(G2072), .A2(G2078), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n442), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  INV_X1    g260(.A(new_n679), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(KEYINPUT17), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(new_n683), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT17), .B1(new_n679), .B2(new_n683), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(new_n681), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n689), .B(new_n691), .C1(new_n686), .C2(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G2096), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n685), .A2(new_n692), .A3(new_n642), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2100), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1971), .B(G1976), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT19), .ZN(new_n705));
  XOR2_X1   g280(.A(G1956), .B(G2474), .Z(new_n706));
  XOR2_X1   g281(.A(G1961), .B(G1966), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(KEYINPUT84), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(KEYINPUT84), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n706), .A2(new_n707), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(new_n708), .ZN(new_n715));
  MUX2_X1   g290(.A(new_n715), .B(new_n714), .S(new_n705), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n712), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1981), .B(G1986), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n703), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n726), .A2(new_n702), .A3(new_n722), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(G229));
  NOR2_X1   g304(.A1(G16), .A2(G22), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G166), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT90), .B(G1971), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  OR2_X1    g309(.A1(G305), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G6), .B2(G16), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT32), .B(G1981), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n735), .B(new_n737), .C1(G6), .C2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n733), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT33), .B(G1976), .Z(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n582), .A2(new_n585), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G16), .ZN(new_n746));
  OR2_X1    g321(.A1(G16), .A2(G23), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n746), .A2(KEYINPUT89), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT89), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n747), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n746), .A2(KEYINPUT89), .A3(new_n747), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(new_n754), .A3(new_n742), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n741), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT91), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n741), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT34), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n758), .A2(KEYINPUT34), .A3(new_n760), .ZN(new_n764));
  NOR2_X1   g339(.A1(G25), .A2(G29), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n640), .A2(G119), .ZN(new_n766));
  NAND2_X1  g341(.A1(G107), .A2(G2105), .ZN(new_n767));
  INV_X1    g342(.A(G95), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G2105), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2104), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G131), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n486), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n766), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n765), .B1(new_n775), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT35), .B(G1991), .Z(new_n777));
  XOR2_X1   g352(.A(new_n776), .B(new_n777), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(KEYINPUT92), .B2(KEYINPUT36), .ZN(new_n779));
  INV_X1    g354(.A(G290), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G16), .B2(G24), .ZN(new_n782));
  INV_X1    g357(.A(G1986), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n779), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n763), .A2(new_n764), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G29), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G33), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n487), .A2(G139), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n464), .A2(new_n466), .A3(G127), .ZN(new_n795));
  INV_X1    g370(.A(G115), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n465), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G2105), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n465), .A2(G2105), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G103), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n794), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n793), .B1(new_n804), .B2(new_n792), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G2072), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n792), .A2(G32), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n487), .A2(G141), .ZN(new_n808));
  NAND3_X1  g383(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT26), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n811), .A2(new_n812), .B1(G105), .B2(new_n799), .ZN(new_n813));
  INV_X1    g388(.A(G129), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n481), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n807), .B1(new_n816), .B2(new_n792), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT27), .B(G1996), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n806), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G29), .A2(G35), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G162), .B2(G29), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT29), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n821), .B1(G2090), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(KEYINPUT24), .A2(G34), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(KEYINPUT24), .A2(G34), .ZN(new_n828));
  AOI21_X1  g403(.A(G29), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G160), .B2(G29), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(G2084), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT31), .B(G11), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT30), .B(G28), .Z(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G29), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n641), .B2(G29), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(G2084), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G1966), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n734), .A2(G21), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G286), .B2(G16), .ZN(new_n840));
  AOI211_X1 g415(.A(new_n831), .B(new_n837), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(G5), .A2(G16), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT94), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G301), .B2(new_n734), .ZN(new_n844));
  INV_X1    g419(.A(G1961), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n840), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n846), .B1(G1966), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n825), .A2(new_n841), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n824), .A2(G2090), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(KEYINPUT96), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n792), .A2(G26), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT28), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n487), .A2(G140), .ZN(new_n855));
  INV_X1    g430(.A(G128), .ZN(new_n856));
  AND2_X1   g431(.A1(G116), .A2(G2105), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G104), .B2(new_n462), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n481), .A2(new_n856), .B1(new_n465), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n854), .B1(new_n860), .B2(new_n792), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G2067), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n845), .B2(new_n844), .ZN(new_n863));
  NOR2_X1   g438(.A1(G27), .A2(G29), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G164), .B2(G29), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT95), .B(G2078), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n852), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n625), .A2(G16), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(G4), .B2(G16), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT93), .B(G1348), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(G16), .A2(G19), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n559), .B2(G16), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(G1341), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n870), .A2(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n734), .A2(G20), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT23), .ZN(new_n878));
  INV_X1    g453(.A(G299), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n734), .ZN(new_n880));
  INV_X1    g455(.A(G1956), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n882), .ZN(new_n883));
  NOR4_X1   g458(.A1(new_n849), .A2(new_n851), .A3(new_n868), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n791), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n786), .B1(new_n761), .B2(new_n762), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n790), .B1(new_n886), .B2(new_n764), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(G311));
  NAND3_X1  g463(.A1(new_n763), .A2(new_n764), .A3(new_n787), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n788), .A3(new_n789), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n791), .A3(new_n884), .ZN(G150));
  AOI22_X1  g466(.A1(G93), .A2(new_n520), .B1(new_n615), .B2(G55), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n531), .A2(G67), .A3(new_n532), .ZN(new_n893));
  NAND2_X1  g468(.A1(G80), .A2(G543), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n503), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G860), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT37), .Z(new_n899));
  NOR2_X1   g474(.A1(new_n620), .A2(new_n626), .ZN(new_n900));
  INV_X1    g475(.A(G93), .ZN(new_n901));
  INV_X1    g476(.A(G55), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n544), .A2(new_n901), .B1(new_n546), .B2(new_n902), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n552), .A2(new_n558), .B1(new_n903), .B2(new_n895), .ZN(new_n904));
  AOI22_X1  g479(.A1(G81), .A2(new_n520), .B1(new_n615), .B2(G43), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n531), .A2(G56), .A3(new_n532), .ZN(new_n906));
  INV_X1    g481(.A(new_n557), .ZN(new_n907));
  OAI21_X1  g482(.A(G651), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n905), .A2(new_n892), .A3(new_n908), .A4(new_n896), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n900), .B(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(KEYINPUT39), .ZN(new_n915));
  INV_X1    g490(.A(G860), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n914), .B2(KEYINPUT39), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n899), .B1(new_n915), .B2(new_n917), .ZN(G145));
  OR3_X1    g493(.A1(new_n462), .A2(KEYINPUT98), .A3(G118), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT98), .B1(new_n462), .B2(G118), .ZN(new_n920));
  OR2_X1    g495(.A1(G106), .A2(G2105), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n919), .A2(G2104), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G130), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n481), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(G142), .B2(new_n487), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n766), .B2(new_n774), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n775), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n647), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(new_n647), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n804), .A2(new_n816), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n860), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n490), .A2(new_n491), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n462), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n493), .A2(new_n494), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G2105), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n939), .A3(new_n498), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n860), .A2(G164), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n804), .A2(new_n816), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n934), .A2(new_n941), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n934), .A2(new_n943), .B1(new_n941), .B2(new_n942), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n929), .B(new_n932), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n932), .A2(new_n929), .ZN(new_n948));
  INV_X1    g523(.A(new_n946), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(G162), .B(new_n479), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(new_n641), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT99), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT99), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n945), .B2(new_n946), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n949), .A2(KEYINPUT100), .A3(new_n944), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n948), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n962), .A2(KEYINPUT101), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT101), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n945), .A2(new_n946), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n953), .B1(new_n965), .B2(new_n948), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n958), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n958), .B2(new_n967), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(G395));
  NOR2_X1   g547(.A1(new_n897), .A2(G868), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n628), .A2(new_n910), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n628), .A2(new_n910), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n977));
  AND3_X1   g552(.A1(new_n612), .A2(new_n879), .A3(new_n619), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n879), .B1(new_n612), .B2(new_n619), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n620), .A2(G299), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n612), .A2(new_n879), .A3(new_n619), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(KEYINPUT41), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n974), .B(new_n975), .C1(new_n979), .C2(new_n978), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G305), .A2(G303), .ZN(new_n988));
  NAND4_X1  g563(.A1(G166), .A2(new_n592), .A3(new_n594), .A4(new_n598), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(new_n744), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n602), .A2(new_n603), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT79), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n604), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n745), .B1(new_n995), .B2(new_n601), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n990), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G290), .A2(new_n744), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n745), .A3(new_n601), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n988), .A4(new_n989), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(KEYINPUT42), .A3(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n987), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n985), .A2(new_n1003), .A3(new_n986), .A4(new_n1004), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n973), .B1(new_n1008), .B2(G868), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(G295));
  XNOR2_X1  g586(.A(new_n1009), .B(KEYINPUT105), .ZN(G331));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n1013));
  INV_X1    g588(.A(new_n977), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n981), .A2(new_n982), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT41), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n978), .B2(new_n979), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n529), .A2(new_n534), .A3(new_n536), .ZN(new_n1018));
  AOI22_X1  g593(.A1(G90), .A2(new_n520), .B1(new_n615), .B2(G52), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n525), .A4(new_n542), .ZN(new_n1020));
  OAI21_X1  g595(.A(G286), .B1(new_n543), .B2(new_n548), .ZN(new_n1021));
  AND4_X1   g596(.A1(new_n904), .A2(new_n909), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n904), .A2(new_n909), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1015), .B(new_n1017), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n910), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n904), .A2(new_n909), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(new_n981), .A3(new_n982), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1001), .A2(KEYINPUT106), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n997), .A2(new_n1031), .A3(new_n1000), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n980), .B(new_n983), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(new_n1001), .A3(new_n1028), .ZN(new_n1035));
  INV_X1    g610(.A(G37), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1013), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1028), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(KEYINPUT43), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT107), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1038), .A2(new_n1042), .A3(new_n1046), .A4(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1039), .A2(new_n1013), .A3(new_n1041), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT108), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1039), .A2(new_n1051), .A3(new_n1013), .A4(new_n1041), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT43), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1050), .A2(KEYINPUT44), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1054), .ZN(G397));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(G164), .B2(G1384), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n467), .A2(new_n468), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G2105), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n470), .B(KEYINPUT69), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n478), .A2(new_n1059), .A3(G40), .A4(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1996), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(KEYINPUT46), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT46), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1062), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n860), .B(G2067), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1069), .A2(new_n816), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1066), .B(new_n1067), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT47), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(KEYINPUT47), .ZN(new_n1074));
  INV_X1    g649(.A(new_n816), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G1996), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1065), .A2(KEYINPUT109), .A3(new_n816), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT109), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1064), .B2(new_n1075), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1077), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n775), .B(new_n777), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1062), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n780), .A2(new_n783), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(new_n1068), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT48), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1073), .A2(new_n1074), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n775), .A2(new_n777), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1089), .B(KEYINPUT125), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n935), .A2(G2067), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1068), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT126), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1087), .A2(new_n1084), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1074), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1072), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1094), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  INV_X1    g678(.A(G1384), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n940), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1061), .B1(new_n1105), .B2(new_n1056), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n940), .A2(KEYINPUT45), .A3(new_n1104), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1971), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n940), .A2(KEYINPUT50), .A3(new_n1104), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1061), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G2090), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1103), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(G303), .A2(G8), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT55), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT63), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1107), .A2(KEYINPUT114), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n940), .A2(new_n1126), .A3(KEYINPUT45), .A4(new_n1104), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1106), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n838), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT115), .B(G2084), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1114), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1103), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G168), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1121), .B1(new_n1124), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1061), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(new_n1104), .A3(new_n940), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G8), .ZN(new_n1137));
  INV_X1    g712(.A(G1976), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n744), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT52), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT111), .ZN(new_n1141));
  INV_X1    g716(.A(G1981), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n592), .A2(new_n1142), .A3(new_n594), .A4(new_n598), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n544), .A2(new_n591), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n597), .A2(G651), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n507), .A2(G48), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(G1981), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1143), .A2(KEYINPUT49), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT49), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1137), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n587), .A2(new_n1138), .A3(new_n588), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT52), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1151), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1134), .A2(new_n1141), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1158), .A2(KEYINPUT63), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT112), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n589), .A2(new_n1160), .A3(new_n1138), .ZN(new_n1161));
  INV_X1    g736(.A(new_n588), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1138), .B1(new_n1162), .B2(new_n586), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT112), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1143), .B1(new_n1165), .B2(new_n1151), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT113), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1137), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT113), .B(new_n1143), .C1(new_n1165), .C2(new_n1151), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1159), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1121), .A2(G168), .A3(new_n1132), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1119), .B1(new_n1172), .B2(new_n1103), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n1141), .A3(new_n1156), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1174), .B2(new_n1122), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1158), .A2(KEYINPUT63), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1157), .B(new_n1170), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G286), .A2(G8), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT123), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT51), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1181));
  OAI211_X1 g756(.A(G8), .B(new_n1180), .C1(new_n1181), .C2(G286), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1180), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1128), .A2(new_n838), .B1(new_n1114), .B2(new_n1130), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1178), .B(new_n1183), .C1(new_n1184), .C2(new_n1103), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1132), .A2(G286), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT62), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1182), .A2(new_n1185), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(G2078), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1106), .A2(new_n1191), .A3(new_n1107), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT53), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n495), .A2(new_n499), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1111), .B(G1384), .C1(new_n1194), .C2(new_n937), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT50), .B1(new_n940), .B2(new_n1104), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1135), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1192), .A2(new_n1193), .B1(new_n1197), .B2(new_n845), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1191), .A2(KEYINPUT53), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1128), .B2(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1200), .A2(G171), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1188), .A2(new_n1190), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1197), .A2(new_n881), .ZN(new_n1203));
  XNOR2_X1  g778(.A(KEYINPUT56), .B(G2072), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1057), .A2(new_n1135), .A3(new_n1107), .A4(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT119), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1106), .A2(KEYINPUT119), .A3(new_n1107), .A4(new_n1204), .ZN(new_n1208));
  AOI21_X1  g783(.A(KEYINPUT57), .B1(new_n572), .B2(KEYINPUT118), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(G299), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1203), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(new_n871), .ZN(new_n1213));
  OAI22_X1  g788(.A1(new_n1114), .A2(new_n1213), .B1(G2067), .B2(new_n1136), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n625), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1203), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1210), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1212), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1214), .A2(KEYINPUT60), .A3(new_n625), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n620), .B(KEYINPUT60), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1136), .A2(G2067), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1222), .B1(new_n1197), .B2(new_n871), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT121), .ZN(new_n1225));
  NOR3_X1   g800(.A1(G164), .A2(G1384), .A3(new_n1061), .ZN(new_n1226));
  XNOR2_X1  g801(.A(KEYINPUT58), .B(G1341), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT120), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1225), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g804(.A1(new_n1057), .A2(new_n1063), .A3(new_n1107), .A4(new_n1135), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1228), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1136), .A2(KEYINPUT121), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT59), .ZN(new_n1234));
  AND3_X1   g809(.A1(new_n1233), .A2(new_n1234), .A3(new_n559), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1234), .B1(new_n1233), .B2(new_n559), .ZN(new_n1236));
  OAI211_X1 g811(.A(new_n1220), .B(new_n1224), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g812(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1211), .ZN(new_n1238));
  NOR2_X1   g813(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1212), .A2(KEYINPUT122), .ZN(new_n1240));
  INV_X1    g815(.A(KEYINPUT122), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1211), .A2(new_n1241), .ZN(new_n1242));
  NAND4_X1  g817(.A1(new_n1240), .A2(KEYINPUT61), .A3(new_n1218), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1219), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g819(.A(G171), .B(KEYINPUT54), .Z(new_n1245));
  AOI21_X1  g820(.A(new_n1199), .B1(new_n1135), .B2(KEYINPUT124), .ZN(new_n1246));
  OAI21_X1  g821(.A(new_n1246), .B1(KEYINPUT124), .B2(new_n1135), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1247), .B1(new_n1056), .B2(new_n1105), .ZN(new_n1248));
  AOI21_X1  g823(.A(new_n1245), .B1(new_n1248), .B2(new_n1107), .ZN(new_n1249));
  AOI22_X1  g824(.A1(new_n1249), .A2(new_n1198), .B1(new_n1200), .B2(new_n1245), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1250), .A2(new_n1187), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1202), .B1(new_n1244), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1174), .B1(new_n1120), .B2(new_n1117), .ZN(new_n1253));
  AOI21_X1  g828(.A(new_n1177), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g829(.A(G290), .B(G1986), .ZN(new_n1255));
  AOI21_X1  g830(.A(new_n1084), .B1(new_n1062), .B2(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g831(.A(new_n1256), .B(KEYINPUT110), .ZN(new_n1257));
  OAI21_X1  g832(.A(new_n1102), .B1(new_n1254), .B2(new_n1257), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g833(.A(new_n460), .B1(new_n674), .B2(new_n675), .ZN(new_n1260));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1261));
  AND3_X1   g835(.A1(new_n1260), .A2(new_n697), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g836(.A(new_n1261), .B1(new_n1260), .B2(new_n697), .ZN(new_n1263));
  OAI21_X1  g837(.A(new_n728), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g838(.A(new_n1264), .B1(new_n958), .B2(new_n967), .ZN(new_n1265));
  AND3_X1   g839(.A1(new_n1265), .A2(new_n1038), .A3(new_n1042), .ZN(G308));
  NAND3_X1  g840(.A1(new_n1265), .A2(new_n1038), .A3(new_n1042), .ZN(G225));
endmodule


