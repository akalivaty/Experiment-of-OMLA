//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT24), .B(G110), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n188), .B2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n189), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT81), .ZN(new_n203));
  AND3_X1   g017(.A1(KEYINPUT80), .A2(G125), .A3(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(G140), .B1(KEYINPUT80), .B2(G125), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n203), .B(KEYINPUT16), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT80), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(KEYINPUT80), .A2(G125), .A3(G140), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n209), .A3(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT81), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n206), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n202), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n196), .A2(new_n189), .A3(new_n197), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G110), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n192), .B2(new_n193), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n206), .B(new_n218), .C1(new_n212), .C2(new_n214), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n216), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(KEYINPUT83), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n202), .A2(new_n220), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(new_n226), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(G953), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n235), .B(KEYINPUT84), .Z(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n221), .A2(new_n227), .A3(new_n235), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n187), .B1(new_n239), .B2(G902), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT25), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G217), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G234), .B2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(G902), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n237), .A2(new_n238), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G469), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G140), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n233), .A2(G227), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT86), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n218), .A2(KEYINPUT66), .A3(G143), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(G146), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n259), .A2(new_n262), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n218), .A2(G143), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n190), .B1(new_n265), .B2(KEYINPUT1), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT3), .B1(new_n268), .B2(G107), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g084(.A(G107), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G104), .ZN(new_n272));
  INV_X1    g086(.A(G101), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(G107), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n269), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n268), .A2(G107), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n271), .A2(G104), .ZN(new_n277));
  OAI21_X1  g091(.A(G101), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n267), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(new_n279), .A3(KEYINPUT85), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT10), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n218), .A2(KEYINPUT64), .A3(G143), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT64), .B1(new_n218), .B2(G143), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n265), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n285), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n265), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n258), .A2(G146), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT64), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT65), .A3(new_n291), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n264), .A2(new_n289), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n269), .A2(new_n272), .A3(new_n274), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G101), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT4), .A3(new_n275), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n304), .A3(G101), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n266), .B1(new_n294), .B2(new_n296), .ZN(new_n307));
  INV_X1    g121(.A(new_n263), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n275), .A2(new_n278), .A3(KEYINPUT10), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n300), .A2(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n256), .B1(new_n284), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n309), .A2(new_n310), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n293), .A2(new_n298), .A3(new_n299), .ZN(new_n314));
  INV_X1    g128(.A(new_n306), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT10), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n267), .A2(new_n279), .A3(KEYINPUT85), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT85), .B1(new_n267), .B2(new_n279), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(KEYINPUT86), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT11), .ZN(new_n323));
  INV_X1    g137(.A(G134), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(G137), .ZN(new_n325));
  INV_X1    g139(.A(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT11), .A3(G134), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(G134), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n322), .B1(new_n330), .B2(new_n323), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n327), .A2(new_n328), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n323), .B1(new_n324), .B2(G137), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT67), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n336), .A4(new_n325), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n312), .A2(new_n321), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n332), .A2(new_n337), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n316), .A2(new_n340), .A3(new_n320), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n255), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n255), .ZN(new_n343));
  INV_X1    g157(.A(new_n279), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n309), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n318), .B2(new_n319), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n346), .A2(KEYINPUT12), .A3(new_n338), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT12), .B1(new_n346), .B2(new_n338), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n251), .B(new_n241), .C1(new_n342), .C2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n341), .B1(new_n347), .B2(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n254), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n284), .A2(new_n311), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n254), .B1(new_n355), .B2(new_n340), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n339), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(G469), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n251), .A2(new_n241), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT9), .B(G234), .ZN(new_n362));
  OAI21_X1  g176(.A(G221), .B1(new_n362), .B2(G902), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G214), .B1(G237), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n233), .A2(G224), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT7), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G125), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n371), .B(new_n263), .C1(new_n288), .C2(new_n266), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT89), .ZN(new_n373));
  INV_X1    g187(.A(new_n266), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n297), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n371), .A4(new_n263), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(KEYINPUT92), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n300), .A2(G125), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(new_n377), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n370), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n188), .A2(G116), .ZN(new_n385));
  INV_X1    g199(.A(G116), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G119), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT2), .B(G113), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT71), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G113), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(KEYINPUT2), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(KEYINPUT2), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n385), .B(new_n387), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(new_n389), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT71), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n303), .A2(new_n391), .A3(new_n397), .A4(new_n305), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n385), .A2(new_n387), .A3(KEYINPUT5), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(G113), .C1(KEYINPUT5), .C2(new_n385), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n279), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G122), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n395), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n344), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n401), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT91), .B(KEYINPUT8), .Z(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n379), .A2(new_n381), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n369), .B1(new_n368), .B2(KEYINPUT93), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(KEYINPUT93), .B2(new_n368), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n403), .B(new_n409), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n241), .B1(new_n384), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n398), .A2(new_n401), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n402), .B(KEYINPUT87), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT88), .ZN(new_n420));
  INV_X1    g234(.A(new_n418), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n398), .B2(new_n401), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n417), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n418), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n403), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n410), .A2(new_n368), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n379), .A2(new_n381), .A3(new_n367), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n425), .A2(KEYINPUT90), .A3(new_n427), .A4(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n403), .A2(KEYINPUT6), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n420), .A2(new_n424), .B1(new_n433), .B2(new_n426), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT90), .B1(new_n434), .B2(new_n430), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n415), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT90), .ZN(new_n440));
  AND4_X1   g254(.A1(new_n423), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n423), .B1(new_n422), .B2(new_n417), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n427), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n428), .A2(new_n429), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n431), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n437), .A3(new_n415), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n366), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n364), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n268), .ZN(new_n451));
  NOR2_X1   g265(.A1(G237), .A2(G953), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G214), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n258), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT18), .A3(G131), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n453), .A2(new_n258), .ZN(new_n456));
  AOI21_X1  g270(.A(G143), .B1(new_n452), .B2(G214), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT18), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n334), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n204), .A2(new_n205), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n219), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT17), .B(G131), .C1(new_n456), .C2(new_n457), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n216), .A2(new_n225), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n216), .A2(KEYINPUT95), .A3(new_n225), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n454), .A2(G131), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n458), .A2(new_n334), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n451), .B(new_n464), .C1(new_n468), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT96), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n466), .A2(new_n467), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n473), .A3(new_n469), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n451), .A4(new_n464), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n470), .A2(new_n471), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT19), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n204), .A2(new_n205), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n485), .B2(new_n217), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n218), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT94), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n484), .A2(new_n216), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n464), .ZN(new_n491));
  INV_X1    g305(.A(new_n451), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n481), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n495));
  NOR2_X1   g309(.A1(G475), .A2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n476), .A2(new_n480), .B1(new_n492), .B2(new_n491), .ZN(new_n498));
  INV_X1    g312(.A(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT20), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n190), .A2(G143), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n258), .A2(G128), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n190), .A2(G143), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT97), .B1(new_n506), .B2(KEYINPUT13), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT97), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n508), .A3(new_n504), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT98), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(G134), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT98), .B1(new_n510), .B2(new_n324), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G116), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n271), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n503), .A2(new_n502), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n324), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n518), .B(new_n324), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n271), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n386), .A2(KEYINPUT14), .A3(G122), .ZN(new_n525));
  INV_X1    g339(.A(new_n516), .ZN(new_n526));
  OAI211_X1 g340(.A(G107), .B(new_n525), .C1(new_n526), .C2(KEYINPUT14), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n362), .A2(new_n244), .A3(G953), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n520), .B1(new_n513), .B2(new_n514), .ZN(new_n532));
  INV_X1    g346(.A(new_n528), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n241), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT99), .B1(new_n535), .B2(new_n241), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n541), .B(G902), .C1(new_n530), .C2(new_n534), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n539), .B1(new_n543), .B2(new_n538), .ZN(new_n544));
  NAND2_X1  g358(.A1(G234), .A2(G237), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(G952), .A3(new_n233), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n545), .A2(G902), .A3(G953), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT21), .B(G898), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n451), .B1(new_n478), .B2(new_n464), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n476), .B2(new_n480), .ZN(new_n552));
  OAI21_X1  g366(.A(G475), .B1(new_n552), .B2(G902), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n501), .A2(new_n544), .A3(new_n550), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n449), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT68), .B1(new_n300), .B2(new_n340), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n330), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n326), .A2(KEYINPUT69), .A3(G134), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n328), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G131), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n337), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT70), .ZN(new_n563));
  INV_X1    g377(.A(new_n309), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n337), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n297), .A2(new_n291), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n568), .A2(new_n285), .B1(new_n264), .B2(new_n289), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT68), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n298), .A4(new_n338), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n556), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n337), .B(new_n561), .C1(new_n307), .C2(new_n308), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT30), .B(new_n575), .C1(new_n300), .C2(new_n340), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n397), .A2(new_n391), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n577), .B(new_n575), .C1(new_n300), .C2(new_n340), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT72), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n452), .A2(G210), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT27), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT26), .B(G101), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n569), .A2(new_n298), .A3(new_n338), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT72), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n577), .A4(new_n575), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n583), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT31), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT74), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n581), .A2(new_n591), .A3(KEYINPUT74), .A4(new_n592), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n579), .B1(new_n573), .B2(new_n572), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n583), .A2(new_n590), .A3(new_n587), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT31), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(KEYINPUT73), .B(KEYINPUT31), .C1(new_n598), .C2(new_n599), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT28), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n582), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n572), .A2(new_n578), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n578), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n583), .A2(new_n590), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT75), .B(KEYINPUT28), .Z(new_n613));
  AOI21_X1  g427(.A(new_n606), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n597), .B(new_n604), .C1(new_n587), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT77), .ZN(new_n616));
  NOR2_X1   g430(.A1(G472), .A2(G902), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT32), .ZN(new_n620));
  INV_X1    g434(.A(new_n617), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT32), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT79), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n615), .A2(KEYINPUT79), .A3(new_n623), .ZN(new_n627));
  INV_X1    g441(.A(new_n587), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n581), .A2(new_n628), .A3(new_n611), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT29), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g445(.A(KEYINPUT29), .B(new_n606), .C1(new_n612), .C2(new_n613), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n575), .B1(new_n300), .B2(new_n340), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n578), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n583), .A2(new_n590), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT28), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n582), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT78), .B1(new_n582), .B2(new_n605), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT29), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n587), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n631), .B1(new_n632), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(G472), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n626), .A2(new_n627), .A3(new_n644), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n250), .B(new_n555), .C1(new_n620), .C2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G101), .ZN(G3));
  NAND2_X1  g461(.A1(new_n615), .A2(new_n617), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT77), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n597), .A2(new_n604), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n614), .A2(new_n587), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n241), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G472), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n649), .A2(new_n653), .A3(new_n654), .A4(new_n364), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n437), .B1(new_n446), .B2(new_n415), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n438), .B(new_n414), .C1(new_n445), .C2(new_n431), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n550), .B(new_n365), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n499), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n553), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n532), .B2(new_n533), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n663), .A2(KEYINPUT33), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n535), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(G478), .A3(new_n241), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n543), .A2(new_n537), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n655), .A2(new_n250), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT101), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n615), .B2(new_n241), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n618), .A2(new_n619), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n661), .ZN(new_n678));
  INV_X1    g492(.A(new_n544), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n658), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n677), .A2(new_n250), .A3(new_n681), .A4(new_n364), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT102), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT35), .B(G107), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  OAI21_X1  g499(.A(new_n365), .B1(new_n656), .B2(new_n657), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n228), .A2(new_n231), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n243), .A2(new_n245), .B1(new_n247), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n686), .A2(new_n554), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n655), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n547), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n546), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n680), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n690), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n364), .A2(new_n448), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n700), .B(new_n703), .C1(new_n620), .C2(new_n645), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  XNOR2_X1  g519(.A(new_n698), .B(KEYINPUT39), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n364), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT40), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n581), .A2(new_n611), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n628), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n241), .B1(new_n635), .B2(new_n587), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n626), .A2(new_n627), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n620), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n656), .A2(new_n657), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n544), .A2(new_n366), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(new_n661), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n690), .ZN(new_n719));
  OR4_X1    g533(.A1(new_n708), .A2(new_n714), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  NAND3_X1  g535(.A1(new_n661), .A2(new_n668), .A3(new_n698), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n703), .B(new_n723), .C1(new_n620), .C2(new_n645), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT103), .B(G146), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G48));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n342), .A2(new_n351), .ZN(new_n728));
  OAI21_X1  g542(.A(G469), .B1(new_n728), .B2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n363), .A3(new_n352), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n250), .B(new_n731), .C1(new_n620), .C2(new_n645), .ZN(new_n732));
  INV_X1    g546(.A(new_n670), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n727), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n615), .A2(KEYINPUT79), .A3(new_n623), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n614), .A2(new_n630), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n587), .A3(new_n641), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n675), .B1(new_n737), .B2(new_n631), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT79), .B1(new_n615), .B2(new_n623), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n649), .A2(new_n622), .A3(new_n654), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n249), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT104), .A3(new_n670), .A4(new_n731), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n734), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NOR2_X1   g560(.A1(new_n735), .A2(new_n739), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n741), .A2(new_n747), .A3(new_n644), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n250), .A3(new_n681), .A4(new_n731), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  NOR4_X1   g564(.A1(new_n686), .A2(new_n730), .A3(new_n554), .A4(new_n690), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n620), .B2(new_n645), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT105), .B(G119), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G21));
  INV_X1    g568(.A(new_n715), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n550), .A2(new_n718), .A3(new_n755), .A4(new_n731), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n640), .A2(new_n628), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n600), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n621), .B1(new_n758), .B2(new_n597), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n652), .B2(G472), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n760), .B2(new_n250), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n676), .A2(new_n762), .A3(new_n249), .A4(new_n759), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n756), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n701), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n686), .A2(new_n730), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n723), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT107), .B(G125), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n358), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n354), .A2(new_n357), .A3(KEYINPUT108), .A4(G469), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n352), .A3(new_n360), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n715), .A2(new_n365), .A3(new_n363), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n722), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n250), .C1(new_n620), .C2(new_n645), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n644), .A2(new_n624), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT32), .B1(new_n615), .B2(new_n617), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n250), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n775), .A2(new_n363), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n656), .A2(new_n657), .A3(new_n366), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n723), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT42), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n778), .A2(KEYINPUT109), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT109), .B1(new_n778), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  NOR3_X1   g603(.A1(new_n776), .A2(new_n680), .A3(new_n699), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n790), .B(new_n250), .C1(new_n620), .C2(new_n645), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n748), .A2(KEYINPUT110), .A3(new_n250), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  AND2_X1   g610(.A1(new_n354), .A2(new_n357), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(KEYINPUT45), .ZN(new_n798));
  OAI21_X1  g612(.A(G469), .B1(new_n797), .B2(KEYINPUT45), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(KEYINPUT46), .A3(new_n360), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n352), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT111), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(KEYINPUT111), .ZN(new_n804));
  INV_X1    g618(.A(new_n800), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n359), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n803), .B(new_n804), .C1(KEYINPUT46), .C2(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n807), .A2(new_n363), .A3(new_n706), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n677), .A2(new_n690), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n678), .A2(new_n668), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(KEYINPUT44), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n809), .A2(new_n812), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT44), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n808), .A2(new_n783), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  INV_X1    g631(.A(new_n783), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n748), .A2(new_n250), .A3(new_n722), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n807), .A2(KEYINPUT47), .A3(new_n363), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT47), .B1(new_n807), .B2(new_n363), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  NAND3_X1  g638(.A1(new_n250), .A2(new_n365), .A3(new_n363), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n729), .A2(new_n352), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n825), .A2(new_n827), .A3(new_n810), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n714), .A2(new_n829), .A3(new_n716), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n702), .B1(new_n740), .B2(new_n741), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n769), .B1(new_n832), .B2(new_n700), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n718), .A2(new_n755), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n775), .A2(new_n690), .A3(new_n363), .A4(new_n698), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n620), .B2(new_n713), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n833), .A2(new_n834), .A3(new_n724), .A4(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n661), .A2(new_n679), .A3(new_n699), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n840), .A2(new_n364), .A3(new_n783), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n620), .B2(new_n645), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n760), .A2(new_n723), .A3(new_n783), .A4(new_n782), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n793), .A2(new_n794), .B1(new_n844), .B2(new_n701), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n766), .A2(new_n768), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n704), .A2(new_n724), .A3(new_n846), .A4(new_n838), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT52), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n788), .A2(new_n839), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n764), .A2(new_n682), .A3(new_n692), .A4(new_n752), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n748), .A2(new_n250), .A3(new_n681), .A4(new_n731), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT112), .B1(new_n658), .B2(new_n669), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n501), .A2(new_n553), .B1(new_n666), .B2(new_n667), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n448), .A2(new_n854), .A3(new_n855), .A4(new_n550), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n655), .A3(new_n250), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT113), .B1(new_n858), .B2(new_n646), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(KEYINPUT113), .A3(new_n646), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n852), .A2(new_n744), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n831), .B1(new_n849), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n839), .A2(new_n848), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n704), .A2(new_n846), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n778), .A2(KEYINPUT53), .A3(new_n785), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n844), .A2(new_n701), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n795), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n748), .A2(new_n751), .B1(new_n655), .B2(new_n691), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n749), .A3(new_n682), .A4(new_n764), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n858), .A2(KEYINPUT113), .A3(new_n646), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n859), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n864), .A2(new_n869), .A3(new_n873), .A4(new_n744), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n863), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n863), .A2(new_n874), .A3(new_n876), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT114), .ZN(new_n879));
  INV_X1    g693(.A(new_n862), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n788), .A2(new_n845), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n866), .A2(new_n831), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n864), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n876), .B1(new_n883), .B2(new_n863), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n887), .B(new_n877), .C1(new_n879), .C2(new_n884), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n818), .A2(new_n730), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n250), .A3(new_n546), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(new_n620), .A3(new_n713), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n661), .A2(new_n668), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n812), .A2(new_n546), .A3(new_n889), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n766), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n716), .A2(new_n366), .A3(new_n731), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT117), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n812), .A2(new_n546), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n761), .A2(new_n763), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT50), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(KEYINPUT50), .A3(new_n908), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n903), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n906), .A2(new_n907), .A3(new_n818), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n807), .A2(new_n363), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT47), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(KEYINPUT116), .A3(new_n820), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n826), .A2(new_n363), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT116), .B1(new_n917), .B2(new_n820), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT51), .B1(new_n913), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n820), .A3(new_n919), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n914), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n901), .A2(new_n912), .A3(new_n925), .A4(KEYINPUT51), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n908), .A2(new_n767), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(G952), .A3(new_n233), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n902), .A2(new_n781), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT48), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n928), .B(new_n930), .C1(new_n855), .C2(new_n894), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n886), .A2(new_n888), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n886), .A2(new_n933), .A3(KEYINPUT120), .A4(new_n888), .ZN(new_n937));
  INV_X1    g751(.A(G952), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n233), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n830), .B1(new_n936), .B2(new_n940), .ZN(G75));
  AOI21_X1  g755(.A(new_n241), .B1(new_n863), .B2(new_n874), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT56), .B1(new_n942), .B2(G210), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n443), .B(new_n430), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n943), .A2(new_n945), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n233), .A2(G952), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(G51));
  NAND2_X1  g763(.A1(new_n863), .A2(new_n874), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT54), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n878), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n359), .B(KEYINPUT57), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n728), .B1(new_n954), .B2(KEYINPUT121), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(KEYINPUT121), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n942), .A2(new_n805), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n948), .B1(new_n956), .B2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n942), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n959), .A2(KEYINPUT122), .A3(new_n498), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT122), .B1(new_n959), .B2(new_n498), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n948), .B1(new_n959), .B2(new_n498), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(new_n886), .A2(new_n888), .ZN(new_n964));
  XOR2_X1   g778(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n965));
  NOR2_X1   g779(.A1(new_n537), .A2(new_n241), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n665), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n952), .A2(new_n665), .A3(new_n967), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n948), .A3(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n863), .B2(new_n874), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n948), .B1(new_n973), .B2(new_n689), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n239), .B(KEYINPUT124), .Z(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT61), .Z(G66));
  INV_X1    g791(.A(new_n548), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n233), .B1(new_n978), .B2(G224), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n862), .B2(new_n233), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n443), .B1(G898), .B2(new_n233), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G69));
  NAND2_X1  g796(.A1(new_n574), .A2(new_n576), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT125), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(new_n487), .Z(new_n985));
  NOR2_X1   g799(.A1(new_n985), .A2(G953), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n833), .A2(new_n724), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT126), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n720), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n823), .A2(new_n816), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n818), .B(new_n707), .C1(new_n669), .C2(new_n680), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n742), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n989), .A2(new_n990), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n986), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(G900), .A2(G953), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n781), .A2(new_n835), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n808), .A2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n1001), .A2(new_n788), .A3(new_n795), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(new_n816), .A3(new_n823), .A4(new_n988), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n999), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n985), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n233), .B1(G227), .B2(G900), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(G72));
  INV_X1    g822(.A(new_n710), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n991), .A2(new_n994), .A3(new_n880), .A4(new_n996), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1003), .B2(new_n862), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n629), .B(KEYINPUT127), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n629), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1009), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n883), .B2(new_n863), .ZN(new_n1019));
  NOR4_X1   g833(.A1(new_n1013), .A2(new_n1016), .A3(new_n948), .A4(new_n1019), .ZN(G57));
endmodule


