//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT85), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT77), .B(G162gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G155gat), .ZN(new_n210));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT78), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n216), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(G155gat), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n219), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n208), .A2(KEYINPUT75), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  AND4_X1   g028(.A1(new_n211), .A2(new_n227), .A3(new_n229), .A4(new_n212), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT74), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G155gat), .B2(G162gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n233), .A3(new_n213), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n226), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n233), .A2(new_n213), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n211), .A2(new_n227), .A3(new_n229), .A4(new_n212), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT76), .A4(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n225), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n224), .A2(new_n217), .B1(new_n235), .B2(new_n238), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G113gat), .B2(G120gat), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(G113gat), .B2(G120gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  INV_X1    g050(.A(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n251), .B(KEYINPUT67), .C1(new_n254), .C2(new_n247), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT68), .B(G113gat), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n256), .A2(new_n253), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n251), .A2(new_n247), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n250), .A2(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n241), .A2(new_n244), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n225), .A3(new_n239), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n240), .A2(new_n260), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n262), .ZN(new_n271));
  INV_X1    g070(.A(new_n268), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n240), .A2(new_n260), .A3(KEYINPUT79), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n267), .A2(new_n268), .B1(new_n274), .B2(KEYINPUT5), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n262), .A2(new_n263), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT4), .B1(new_n242), .B2(new_n259), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n241), .A2(new_n244), .A3(new_n260), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n268), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n207), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(KEYINPUT5), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n267), .A2(KEYINPUT5), .A3(new_n268), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT86), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n206), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT40), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT39), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n292), .B(new_n272), .C1(new_n261), .C2(new_n266), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n206), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n272), .B1(new_n261), .B2(new_n266), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n271), .A2(new_n273), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n297), .B(KEYINPUT39), .C1(new_n272), .C2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(KEYINPUT40), .A3(new_n206), .A4(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n288), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G211gat), .B(G218gat), .Z(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G226gat), .ZN(new_n311));
  INV_X1    g110(.A(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n321), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(KEYINPUT64), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n319), .B(new_n320), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n317), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n326), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n327), .B2(new_n326), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n319), .A2(new_n320), .ZN(new_n334));
  INV_X1    g133(.A(new_n318), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n321), .A2(KEYINPUT23), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n323), .A2(KEYINPUT64), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n333), .A2(new_n334), .A3(new_n316), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n335), .A2(KEYINPUT26), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  INV_X1    g143(.A(G169gat), .ZN(new_n345));
  INV_X1    g144(.A(G176gat), .ZN(new_n346));
  AND4_X1   g145(.A1(KEYINPUT66), .A2(new_n344), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT66), .B1(new_n318), .B2(new_n344), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n343), .B(new_n320), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT27), .B(G183gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT28), .B1(new_n352), .B2(new_n327), .ZN(new_n353));
  INV_X1    g152(.A(G183gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT27), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G183gat), .ZN(new_n357));
  AND4_X1   g156(.A1(KEYINPUT28), .A2(new_n355), .A3(new_n357), .A4(new_n327), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n315), .B1(new_n342), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n331), .A2(new_n339), .B1(KEYINPUT65), .B2(KEYINPUT25), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n351), .A2(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(new_n313), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n310), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n360), .A3(new_n313), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n314), .B1(new_n362), .B2(new_n363), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n308), .B(new_n309), .Z(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(KEYINPUT71), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n372), .B(new_n310), .C1(new_n361), .C2(new_n365), .ZN(new_n373));
  XOR2_X1   g172(.A(G8gat), .B(G36gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT72), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n371), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n371), .A2(new_n373), .B1(KEYINPUT30), .B2(new_n378), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n371), .B2(new_n373), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n379), .A2(new_n380), .B1(new_n381), .B2(KEYINPUT30), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n371), .A2(new_n373), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n378), .A2(KEYINPUT30), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n373), .A3(new_n378), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n378), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT84), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n384), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n302), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n310), .B1(new_n244), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n308), .A2(new_n400), .A3(new_n309), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n401), .B(new_n398), .C1(new_n310), .C2(new_n400), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n242), .B1(new_n402), .B2(new_n243), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n310), .B2(new_n398), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n242), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n404), .A2(new_n405), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(KEYINPUT82), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n415), .B2(new_n412), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n408), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n285), .A2(new_n286), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n419), .A2(new_n420), .A3(new_n205), .ZN(new_n421));
  INV_X1    g220(.A(new_n206), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n275), .A2(new_n282), .A3(new_n207), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT86), .B1(new_n285), .B2(new_n286), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT6), .B1(new_n419), .B2(new_n205), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n378), .B1(new_n385), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n366), .A2(new_n370), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT38), .B1(new_n430), .B2(KEYINPUT37), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n390), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT38), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n371), .A2(KEYINPUT37), .A3(new_n373), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n418), .B1(new_n427), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n302), .A2(new_n394), .A3(KEYINPUT87), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n397), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n417), .B(KEYINPUT83), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n419), .A2(new_n205), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n421), .B1(new_n442), .B2(new_n426), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n389), .A2(KEYINPUT73), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT73), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n387), .A2(new_n445), .A3(new_n388), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n392), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT69), .B(G71gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(G99gat), .ZN(new_n451));
  XOR2_X1   g250(.A(G15gat), .B(G43gat), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n342), .A2(new_n260), .A3(new_n360), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n259), .B1(new_n362), .B2(new_n363), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n456), .B2(KEYINPUT70), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n454), .A2(new_n455), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n457), .B(new_n462), .C1(new_n454), .C2(new_n455), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n460), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n458), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n467), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n449), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n458), .A2(KEYINPUT32), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT36), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n448), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n472), .B2(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT88), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n427), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n384), .A2(new_n393), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n418), .A2(KEYINPUT35), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n442), .A2(new_n426), .ZN(new_n490));
  INV_X1    g289(.A(new_n421), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n418), .A2(new_n472), .A3(new_n473), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n444), .A2(new_n392), .A3(new_n446), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n440), .A2(new_n481), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT16), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n498), .B(KEYINPUT93), .C1(new_n499), .C2(G1gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n414), .A2(G15gat), .ZN(new_n501));
  INV_X1    g300(.A(G15gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G22gat), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n501), .B(new_n503), .C1(new_n499), .C2(G1gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(G1gat), .B1(new_n501), .B2(new_n503), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT94), .B(G8gat), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n500), .A2(new_n506), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n504), .B(KEYINPUT92), .C1(G1gat), .C2(new_n498), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n520), .A2(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n519), .ZN(new_n532));
  NAND2_X1  g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n522), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n536), .A3(KEYINPUT15), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n527), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(new_n532), .A3(new_n536), .A4(KEYINPUT15), .ZN(new_n541));
  AOI211_X1 g340(.A(KEYINPUT91), .B(new_n518), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n538), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT15), .B1(new_n532), .B2(new_n536), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT17), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n517), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n539), .A2(new_n541), .B1(new_n510), .B2(new_n515), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n549), .A4(new_n551), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n549), .B(KEYINPUT13), .Z(new_n556));
  NOR2_X1   g355(.A1(new_n516), .A2(new_n545), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n560), .B(new_n556), .C1(new_n557), .C2(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n554), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(G169gat), .B(G197gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT12), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n562), .A4(new_n569), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT96), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n563), .A2(new_n574), .A3(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n545), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT8), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n586), .A2(KEYINPUT100), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT100), .B1(new_n586), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n595), .B(new_n584), .C1(new_n590), .C2(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT101), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n542), .B2(new_n547), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n599), .B2(new_n600), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n580), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n603), .A3(new_n579), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G57gat), .B(G64gat), .Z(new_n611));
  OR2_X1    g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G57gat), .B(G64gat), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n613), .B(new_n612), .C1(new_n618), .C2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT99), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G183gat), .B(G211gat), .Z(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n517), .B1(new_n620), .B2(new_n621), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n634), .B(new_n637), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n632), .B2(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n610), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n617), .A2(new_n619), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n594), .A2(new_n643), .A3(new_n596), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n597), .A2(new_n620), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT10), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n644), .ZN(new_n653));
  INV_X1    g452(.A(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n652), .A2(new_n655), .A3(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n497), .A2(new_n576), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n443), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(new_n394), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n670), .A2(new_n672), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(G8gat), .B2(new_n670), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n675), .B2(new_n669), .ZN(G1325gat));
  NAND3_X1  g475(.A1(new_n666), .A2(new_n502), .A3(new_n485), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n480), .A2(KEYINPUT103), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n480), .A2(KEYINPUT103), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n666), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(new_n681), .B2(new_n502), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n441), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n497), .A2(new_n609), .ZN(new_n686));
  INV_X1    g485(.A(new_n641), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n663), .ZN(new_n688));
  INV_X1    g487(.A(new_n576), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n492), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n497), .B2(new_n609), .ZN(new_n696));
  NAND2_X1  g495(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n448), .A2(new_n480), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n302), .A2(new_n394), .A3(KEYINPUT87), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT87), .B1(new_n302), .B2(new_n394), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n698), .B1(new_n701), .B2(new_n438), .ZN(new_n702));
  AND4_X1   g501(.A1(new_n487), .A2(new_n484), .A3(new_n483), .A4(new_n488), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n703), .A2(new_n486), .B1(KEYINPUT35), .B2(new_n495), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n610), .B(new_n697), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n690), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(new_n443), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n694), .B1(new_n529), .B2(new_n707), .ZN(G1328gat));
  NAND4_X1  g507(.A1(new_n688), .A2(new_n530), .A3(new_n394), .A4(new_n610), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n497), .A2(new_n576), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT46), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n706), .A2(new_n394), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n530), .ZN(G1329gat));
  XOR2_X1   g512(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n714));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n686), .A2(new_n715), .A3(new_n485), .A4(new_n691), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT106), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n706), .B2(new_n680), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n480), .B(new_n690), .C1(new_n696), .C2(new_n705), .ZN(new_n720));
  OAI211_X1 g519(.A(KEYINPUT47), .B(new_n716), .C1(new_n720), .C2(new_n715), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(new_n441), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n692), .A2(KEYINPUT107), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n441), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(G50gat), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n706), .B2(new_n418), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n692), .A2(new_n725), .B1(KEYINPUT107), .B2(KEYINPUT48), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n728), .A2(KEYINPUT48), .B1(new_n730), .B2(new_n731), .ZN(G1331gat));
  NAND3_X1  g531(.A1(new_n642), .A2(new_n576), .A3(new_n663), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n497), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n443), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g535(.A1(new_n497), .A2(new_n487), .A3(new_n733), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  AND2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n737), .B2(new_n738), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n485), .ZN(new_n742));
  AOI21_X1  g541(.A(G71gat), .B1(new_n742), .B2(KEYINPUT108), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(KEYINPUT108), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n734), .A2(G71gat), .A3(new_n680), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n441), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT110), .B(G78gat), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1335gat));
  NOR2_X1   g551(.A1(new_n689), .A2(new_n687), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n610), .B(new_n753), .C1(new_n702), .C2(new_n704), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(KEYINPUT51), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n492), .A2(G85gat), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n755), .A2(new_n663), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n663), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n696), .B2(new_n705), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n443), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(new_n587), .ZN(G1336gat));
  NOR2_X1   g561(.A1(new_n487), .A2(G92gat), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n755), .A2(new_n663), .A3(new_n756), .A4(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n760), .A2(new_n394), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n588), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n768), .B(new_n764), .C1(new_n765), .C2(new_n588), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(new_n485), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(G99gat), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n663), .A3(new_n756), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n760), .A2(new_n680), .ZN(new_n774));
  INV_X1    g573(.A(G99gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(G1338gat));
  NOR2_X1   g575(.A1(new_n417), .A2(G106gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n663), .A3(new_n756), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n760), .B2(new_n441), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n780), .B2(KEYINPUT111), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n782), .B(new_n779), .C1(new_n760), .C2(new_n441), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT53), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n760), .A2(new_n418), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(new_n778), .C1(new_n786), .C2(new_n779), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1339gat));
  NAND2_X1  g587(.A1(new_n651), .A2(new_n650), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT10), .B1(new_n644), .B2(new_n645), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n654), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(KEYINPUT54), .A3(new_n652), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n651), .A2(new_n650), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n649), .A4(new_n648), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n660), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(new_n662), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n791), .A2(KEYINPUT54), .A3(new_n652), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n660), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n573), .A2(new_n797), .A3(new_n575), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n549), .B1(new_n548), .B2(new_n551), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n557), .A2(new_n550), .A3(new_n556), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n568), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n663), .A2(new_n572), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n610), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n801), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n572), .A2(new_n805), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(new_n609), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n641), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n642), .A2(new_n576), .A3(new_n664), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n492), .A2(new_n394), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n493), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n256), .A3(new_n689), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n441), .B1(new_n811), .B2(new_n812), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n814), .A2(new_n485), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n576), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(G1340gat));
  AOI21_X1  g622(.A(new_n253), .B1(new_n820), .B2(new_n663), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT112), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n816), .A2(new_n253), .A3(new_n663), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n816), .A2(new_n828), .A3(new_n687), .ZN(new_n829));
  OAI21_X1  g628(.A(G127gat), .B1(new_n821), .B2(new_n641), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1342gat));
  INV_X1    g630(.A(G134gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n832), .A3(new_n610), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n821), .B2(new_n609), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n680), .A2(new_n417), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n815), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(G141gat), .B1(new_n840), .B2(new_n689), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(KEYINPUT116), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n813), .A2(new_n845), .A3(new_n418), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n814), .A2(new_n480), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n552), .A2(new_n553), .B1(new_n559), .B2(new_n561), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n569), .B1(new_n850), .B2(new_n555), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n799), .B2(new_n800), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n662), .A3(new_n796), .ZN(new_n855));
  INV_X1    g654(.A(new_n575), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n663), .A2(new_n572), .A3(new_n859), .A4(new_n805), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT115), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n573), .A2(new_n797), .A3(new_n575), .A4(new_n854), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n863), .A2(new_n864), .A3(new_n858), .A4(new_n860), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n609), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n810), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n687), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n812), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n441), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n848), .B1(KEYINPUT57), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(G141gat), .A3(new_n689), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n843), .A2(new_n844), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n844), .B1(new_n843), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G148gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n871), .B2(new_n663), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n802), .A2(new_n806), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n609), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n687), .B1(new_n881), .B2(new_n867), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT57), .B(new_n418), .C1(new_n882), .C2(new_n869), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n813), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n418), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n845), .A2(new_n870), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n847), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n847), .A2(new_n888), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n663), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G148gat), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n879), .B1(new_n892), .B2(KEYINPUT59), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n839), .A2(G148gat), .A3(new_n664), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n876), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n894), .ZN(new_n896));
  INV_X1    g695(.A(new_n891), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n885), .A2(new_n886), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n863), .A2(new_n858), .A3(new_n860), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n610), .B1(new_n899), .B2(KEYINPUT115), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n810), .B1(new_n900), .B2(new_n865), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n812), .B1(new_n901), .B2(new_n687), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n441), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n897), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n877), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT119), .B(new_n896), .C1(new_n905), .C2(new_n879), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n895), .A2(new_n906), .ZN(G1345gat));
  INV_X1    g706(.A(G155gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n871), .B2(new_n687), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n839), .A2(G155gat), .A3(new_n641), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n909), .A2(new_n910), .ZN(G1346gat));
  OR3_X1    g710(.A1(new_n839), .A2(new_n209), .A3(new_n609), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n871), .A2(KEYINPUT120), .A3(new_n610), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n209), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT120), .B1(new_n871), .B2(new_n610), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(G1347gat));
  INV_X1    g715(.A(new_n493), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n487), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n443), .B1(new_n811), .B2(new_n812), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n689), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n492), .A2(new_n394), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n771), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n818), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n818), .A2(KEYINPUT122), .A3(new_n924), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n576), .A2(new_n345), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n922), .B1(new_n929), .B2(new_n930), .ZN(G1348gat));
  NAND3_X1  g730(.A1(new_n921), .A2(new_n346), .A3(new_n663), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n929), .A2(new_n663), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n346), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n927), .A2(new_n687), .A3(new_n928), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n927), .A2(new_n937), .A3(new_n687), .A4(new_n928), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(G183gat), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n352), .A3(new_n687), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g740(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n327), .A3(new_n610), .ZN(new_n944));
  INV_X1    g743(.A(new_n929), .ZN(new_n945));
  OAI21_X1  g744(.A(G190gat), .B1(new_n945), .B2(new_n609), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(KEYINPUT61), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  NAND3_X1  g748(.A1(new_n838), .A2(KEYINPUT125), .A3(new_n394), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n418), .B(new_n394), .C1(new_n678), .C2(new_n679), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n953), .A3(new_n920), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n689), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n887), .A2(new_n680), .A3(new_n923), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n689), .A2(G197gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n663), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G204gat), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n664), .A2(G204gat), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n950), .A2(new_n953), .A3(new_n920), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n965));
  XOR2_X1   g764(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n966));
  OAI211_X1 g765(.A(new_n961), .B(new_n965), .C1(new_n964), .C2(new_n966), .ZN(G1353gat));
  NOR2_X1   g766(.A1(new_n680), .A2(new_n923), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n687), .B(new_n968), .C1(new_n898), .C2(new_n903), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n687), .A2(new_n305), .ZN(new_n972));
  OAI22_X1  g771(.A1(new_n970), .A2(new_n971), .B1(new_n954), .B2(new_n972), .ZN(G1354gat));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n306), .A3(new_n610), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n957), .A2(new_n610), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n306), .ZN(G1355gat));
endmodule


