//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n206), .C1(new_n207), .C2(KEYINPUT2), .ZN(new_n208));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT76), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(new_n207), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n203), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT76), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n208), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G113gat), .ZN(new_n224));
  INV_X1    g023(.A(G113gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G120gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT1), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G127gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G134gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G134gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G127gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n233), .A3(KEYINPUT67), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n227), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n233), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n206), .A2(new_n203), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n210), .B2(new_n220), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n213), .B1(new_n212), .B2(new_n207), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n215), .A2(KEYINPUT76), .A3(new_n220), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n236), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n230), .B1(new_n246), .B2(KEYINPUT67), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n247), .B2(new_n227), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT78), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254));
  AOI211_X1 g053(.A(new_n254), .B(new_n251), .C1(new_n239), .C2(new_n249), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n222), .A2(new_n258), .A3(KEYINPUT3), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT77), .B1(new_n244), .B2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n238), .B(new_n257), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT4), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT4), .B1(new_n244), .B2(new_n248), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n265), .A3(new_n251), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n262), .A2(new_n265), .A3(new_n251), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT81), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n271), .A2(new_n276), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n280));
  INV_X1    g079(.A(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n268), .A2(new_n281), .A3(new_n270), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n271), .A2(new_n284), .A3(KEYINPUT6), .A4(new_n276), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n278), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G226gat), .ZN(new_n287));
  INV_X1    g086(.A(G233gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT23), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT24), .ZN(new_n299));
  NOR2_X1   g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n293), .A2(new_n295), .A3(new_n303), .A4(new_n296), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n298), .A2(KEYINPUT24), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(KEYINPUT25), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT24), .A3(new_n298), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n312), .A2(new_n296), .A3(new_n295), .A4(new_n293), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n308), .B1(new_n313), .B2(new_n305), .ZN(new_n314));
  INV_X1    g113(.A(new_n298), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT26), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n296), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n292), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(KEYINPUT65), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT65), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NOR4_X1   g123(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n322), .B2(new_n316), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n315), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT27), .B(G183gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n310), .ZN(new_n332));
  AND2_X1   g131(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n310), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n307), .A2(new_n314), .B1(new_n329), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n290), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n338), .B2(new_n290), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n328), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n342), .A3(new_n298), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n302), .A2(new_n306), .B1(KEYINPUT25), .B2(new_n304), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n293), .A2(new_n295), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(new_n296), .A3(new_n306), .A4(new_n312), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n308), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT73), .A3(new_n289), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(new_n341), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  INV_X1    g151(.A(G211gat), .ZN(new_n353));
  INV_X1    g152(.A(G218gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n351), .A3(new_n355), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT70), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n362), .A3(new_n358), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n361), .A2(KEYINPUT71), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT71), .B1(new_n361), .B2(new_n363), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n307), .A2(new_n314), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n368), .B2(new_n343), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT72), .B1(new_n369), .B2(new_n289), .ZN(new_n370));
  INV_X1    g169(.A(new_n366), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n348), .A2(new_n289), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n290), .C1(new_n338), .C2(KEYINPUT29), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n370), .A2(new_n371), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n367), .B2(new_n375), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(KEYINPUT30), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n376), .A2(KEYINPUT30), .A3(new_n380), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n380), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n202), .B1(new_n286), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n278), .A2(new_n283), .A3(new_n285), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n383), .B2(new_n386), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n398), .A4(new_n392), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT31), .ZN(new_n401));
  XOR2_X1   g200(.A(KEYINPUT83), .B(G50gat), .Z(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n258), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n244), .A2(KEYINPUT77), .A3(new_n260), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n366), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n359), .A2(new_n409), .A3(new_n360), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n410), .B(new_n411), .C1(new_n409), .C2(new_n360), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n244), .B1(new_n412), .B2(new_n260), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n404), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n404), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n361), .A2(new_n411), .A3(new_n363), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n417), .A2(new_n260), .ZN(new_n418));
  OAI221_X1 g217(.A(new_n416), .B1(new_n418), .B2(new_n244), .C1(new_n407), .C2(new_n366), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n414), .B2(new_n419), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n403), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n403), .A2(KEYINPUT85), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(KEYINPUT85), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n396), .A2(new_n399), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n376), .A2(KEYINPUT37), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n350), .A2(new_n371), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n370), .A2(new_n366), .A3(new_n372), .A4(new_n374), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n433), .A2(KEYINPUT37), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n379), .B(new_n431), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n376), .A2(KEYINPUT37), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n379), .B1(new_n437), .B2(new_n432), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n385), .B1(new_n438), .B2(new_n430), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n286), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n262), .A2(KEYINPUT39), .A3(new_n265), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT39), .B1(new_n262), .B2(new_n265), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n252), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n250), .A2(KEYINPUT39), .A3(new_n251), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n281), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n395), .A2(new_n279), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n428), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n440), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n348), .A2(new_n238), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n338), .A2(new_n248), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n455), .B2(KEYINPUT68), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n368), .A2(new_n248), .A3(new_n343), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n248), .B1(new_n368), .B2(new_n343), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n456), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G43gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  AOI21_X1  g268(.A(new_n461), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  AOI211_X1 g270(.A(new_n460), .B(new_n471), .C1(new_n464), .C2(new_n465), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n455), .B1(new_n452), .B2(new_n453), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n469), .B1(new_n476), .B2(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n460), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n466), .A2(new_n461), .A3(new_n469), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n458), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n474), .B1(new_n470), .B2(new_n472), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n473), .A3(new_n479), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n457), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT69), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT36), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n482), .A2(new_n457), .A3(new_n483), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n457), .B1(new_n482), .B2(new_n483), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n429), .A2(new_n451), .A3(new_n487), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n396), .A2(new_n399), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n485), .A2(new_n428), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n286), .A2(new_n395), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(KEYINPUT87), .A3(new_n494), .A4(new_n496), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n423), .A2(new_n427), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(new_n484), .A3(new_n481), .A4(new_n426), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n397), .A2(new_n494), .A3(new_n398), .A4(new_n392), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n493), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT89), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(G29gat), .A3(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  XOR2_X1   g312(.A(G43gat), .B(G50gat), .Z(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n513), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT90), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n515), .A2(new_n516), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n514), .A2(new_n513), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n512), .B2(new_n520), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT91), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT17), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  OR3_X1    g328(.A1(new_n529), .A2(KEYINPUT92), .A3(G1gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT92), .B1(new_n529), .B2(G1gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT93), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT93), .B1(new_n531), .B2(G1gat), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n534), .B(G8gat), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n531), .A2(G1gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n533), .B2(KEYINPUT94), .ZN(new_n539));
  INV_X1    g338(.A(G8gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(new_n540), .C1(KEYINPUT94), .C2(new_n533), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n526), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT18), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n542), .B(new_n545), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n547), .B(KEYINPUT13), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(KEYINPUT18), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n555));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT12), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n549), .A2(new_n560), .A3(new_n553), .A4(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G230gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(new_n288), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n570));
  AOI211_X1 g369(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n570), .B2(KEYINPUT7), .ZN(new_n572));
  INV_X1    g371(.A(G99gat), .ZN(new_n573));
  INV_X1    g372(.A(G106gat), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT8), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT98), .B(G85gat), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n569), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578));
  OAI211_X1 g377(.A(KEYINPUT97), .B(new_n578), .C1(new_n568), .C2(new_n569), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n572), .A2(new_n575), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G99gat), .B(G106gat), .Z(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(KEYINPUT95), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G71gat), .B(G78gat), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n587), .B(new_n588), .C1(KEYINPUT95), .C2(new_n586), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n582), .A2(new_n583), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n593), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n567), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n567), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n595), .B2(new_n598), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n565), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n542), .B1(KEYINPUT21), .B2(new_n594), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G183gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT20), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n615), .B(new_n617), .Z(new_n618));
  NOR2_X1   g417(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n618), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n528), .A2(new_n597), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n584), .A2(new_n545), .ZN(new_n626));
  NAND3_X1  g425(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(KEYINPUT99), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n632), .A2(KEYINPUT100), .ZN(new_n633));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(KEYINPUT100), .ZN(new_n637));
  AND4_X1   g436(.A1(new_n631), .A2(new_n633), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n633), .A2(new_n637), .B1(new_n631), .B2(new_n636), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n506), .A2(new_n611), .A3(new_n624), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n286), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g443(.A1(new_n642), .A2(new_n395), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n648), .B(new_n649), .C1(new_n540), .C2(new_n645), .ZN(G1325gat));
  INV_X1    g449(.A(new_n485), .ZN(new_n651));
  AOI21_X1  g450(.A(G15gat), .B1(new_n642), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n492), .A2(KEYINPUT102), .A3(new_n487), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT102), .B1(new_n492), .B2(new_n487), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n642), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n652), .B1(G15gat), .B2(new_n656), .ZN(G1326gat));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n428), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  INV_X1    g459(.A(new_n640), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n662));
  AOI21_X1  g461(.A(new_n502), .B1(new_n396), .B2(new_n399), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n504), .B(new_n499), .C1(new_n663), .C2(new_n494), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n429), .B(new_n451), .C1(new_n653), .C2(new_n654), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT106), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT106), .B1(new_n664), .B2(new_n665), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n661), .B(new_n662), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n506), .A2(new_n661), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT105), .B1(new_n669), .B2(KEYINPUT44), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n640), .B1(new_n664), .B2(new_n493), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n668), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n610), .B(KEYINPUT103), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n623), .A3(new_n564), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT104), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT108), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n397), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n669), .A2(new_n624), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n611), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n683), .A2(G29gat), .A3(new_n397), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT45), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(G1328gat));
  INV_X1    g485(.A(new_n395), .ZN(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n680), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n683), .A2(G36gat), .A3(new_n687), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(new_n655), .ZN(new_n692));
  OAI21_X1  g491(.A(G43gat), .B1(new_n679), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n683), .A2(G43gat), .A3(new_n485), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(KEYINPUT47), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n680), .A2(new_n692), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n694), .B1(new_n697), .B2(G43gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g498(.A(G50gat), .B1(new_n679), .B2(new_n450), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n683), .A2(G50gat), .A3(new_n450), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n680), .A2(new_n450), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(G50gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n666), .A2(new_n667), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n676), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n661), .A2(new_n564), .A3(new_n623), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n286), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g512(.A(new_n687), .B(new_n710), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1333gat));
  NAND3_X1  g515(.A1(new_n711), .A2(G71gat), .A3(new_n655), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n710), .A2(new_n485), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(G71gat), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n711), .A2(new_n428), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n623), .A2(new_n565), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n664), .B2(new_n665), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n661), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT51), .B1(new_n724), .B2(new_n661), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n610), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n286), .A3(new_n576), .ZN(new_n729));
  INV_X1    g528(.A(new_n610), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n669), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI211_X1 g534(.A(KEYINPUT109), .B(new_n732), .C1(new_n735), .C2(new_n668), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n675), .B2(new_n731), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n397), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n729), .B1(new_n740), .B2(new_n576), .ZN(G1336gat));
  INV_X1    g540(.A(new_n676), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n569), .B(new_n742), .C1(new_n725), .C2(new_n726), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n687), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n395), .B1(new_n736), .B2(new_n738), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(G92gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n732), .B1(new_n735), .B2(new_n668), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n569), .B1(new_n748), .B2(new_n395), .ZN(new_n749));
  NOR4_X1   g548(.A1(new_n749), .A2(new_n744), .A3(KEYINPUT110), .A4(KEYINPUT52), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n675), .A2(new_n395), .A3(new_n731), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(new_n752), .B2(G92gat), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n743), .A2(new_n687), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n746), .A2(new_n747), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(G92gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n747), .A3(new_n754), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n753), .A2(new_n751), .A3(new_n754), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n762), .B(new_n763), .C1(new_n747), .C2(new_n746), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n757), .A2(new_n764), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n739), .B2(new_n692), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n728), .A2(new_n573), .A3(new_n651), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(G1338gat));
  NAND2_X1  g567(.A1(new_n675), .A2(new_n731), .ZN(new_n769));
  OAI21_X1  g568(.A(G106gat), .B1(new_n769), .B2(new_n450), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n727), .A2(new_n574), .A3(new_n428), .A4(new_n742), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n748), .A2(new_n737), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n450), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT112), .B1(new_n776), .B2(new_n574), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n778), .B(G106gat), .C1(new_n739), .C2(new_n450), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n780), .B2(new_n771), .ZN(G1339gat));
  AOI21_X1  g580(.A(new_n547), .B1(new_n544), .B2(new_n546), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n550), .A2(new_n551), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n785), .A2(new_n786), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n559), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n610), .A2(new_n563), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n599), .A2(new_n600), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n602), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n599), .A2(new_n600), .A3(new_n567), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n607), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n601), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT113), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n795), .A2(new_n798), .A3(new_n803), .A4(KEYINPUT55), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n801), .A2(new_n608), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n791), .B1(new_n805), .B2(new_n565), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT116), .B(new_n791), .C1(new_n805), .C2(new_n565), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n640), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n805), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n790), .A2(new_n563), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n811), .B(new_n812), .C1(new_n638), .C2(new_n639), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n624), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n661), .A2(new_n623), .A3(new_n610), .A4(new_n564), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n286), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n687), .A3(new_n496), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n565), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n496), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n687), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n564), .A2(new_n225), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  NAND2_X1  g623(.A1(new_n610), .A2(new_n223), .ZN(new_n825));
  OAI21_X1  g624(.A(G120gat), .B1(new_n818), .B2(new_n676), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n822), .A2(new_n825), .B1(new_n828), .B2(new_n829), .ZN(G1341gat));
  NOR3_X1   g629(.A1(new_n818), .A2(new_n228), .A3(new_n623), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n821), .A2(new_n687), .A3(new_n624), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n228), .ZN(G1342gat));
  NOR2_X1   g632(.A1(new_n640), .A2(new_n395), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n821), .A2(new_n232), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n818), .B2(new_n640), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n838), .A3(new_n232), .A4(new_n834), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(G1343gat));
  OAI21_X1  g639(.A(new_n428), .B1(new_n814), .B2(new_n815), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n655), .A2(new_n397), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n687), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(G141gat), .A3(new_n565), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n791), .A2(KEYINPUT120), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n801), .A2(new_n804), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n799), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(KEYINPUT122), .A2(KEYINPUT55), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n795), .A2(KEYINPUT121), .A3(new_n798), .ZN(new_n857));
  NAND2_X1  g656(.A1(KEYINPUT122), .A2(KEYINPUT55), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n853), .A2(new_n608), .A3(new_n564), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n791), .A2(KEYINPUT120), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n852), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n640), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n624), .B1(new_n863), .B2(new_n813), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n428), .B1(new_n864), .B2(new_n815), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(new_n848), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n841), .A2(KEYINPUT119), .A3(new_n848), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n564), .A3(new_n845), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n847), .B1(new_n869), .B2(G141gat), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT123), .B1(new_n869), .B2(G141gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  AOI221_X4 g672(.A(new_n847), .B1(KEYINPUT123), .B2(new_n873), .C1(new_n869), .C2(G141gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(G1344gat));
  AND2_X1   g674(.A1(new_n868), .A2(new_n845), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n216), .C1(new_n876), .C2(new_n610), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n865), .B2(new_n848), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n848), .B2(new_n841), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n842), .A2(new_n879), .A3(KEYINPUT57), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n610), .A3(new_n845), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n610), .A2(new_n216), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n877), .A2(new_n884), .B1(new_n846), .B2(new_n885), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n846), .A2(new_n623), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT125), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n623), .A2(new_n204), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n888), .A2(new_n204), .B1(new_n876), .B2(new_n889), .ZN(G1346gat));
  NAND2_X1  g689(.A1(new_n876), .A2(new_n661), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n876), .A2(KEYINPUT126), .A3(new_n661), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(G162gat), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n842), .A2(new_n205), .A3(new_n834), .A4(new_n843), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1347gat));
  AND2_X1   g696(.A1(new_n816), .A2(new_n397), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n395), .A3(new_n496), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n565), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(new_n291), .ZN(G1348gat));
  NOR3_X1   g700(.A1(new_n899), .A2(new_n292), .A3(new_n676), .ZN(new_n902));
  INV_X1    g701(.A(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n610), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n292), .B2(new_n904), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n899), .A2(new_n623), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n331), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n309), .B2(new_n906), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G190gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n899), .A2(new_n640), .ZN(new_n912));
  MUX2_X1   g711(.A(new_n910), .B(new_n911), .S(new_n912), .Z(G1351gat));
  NOR2_X1   g712(.A1(new_n655), .A2(new_n286), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n881), .A2(new_n395), .A3(new_n882), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n565), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n692), .A2(new_n395), .A3(new_n428), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n898), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n565), .A2(G197gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  NOR3_X1   g721(.A1(new_n920), .A2(G204gat), .A3(new_n730), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g725(.A(G204gat), .B1(new_n915), .B2(new_n676), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G1353gat));
  INV_X1    g727(.A(new_n920), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n353), .A3(new_n624), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n915), .A2(new_n623), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n932));
  OAI211_X1 g731(.A(KEYINPUT63), .B(G211gat), .C1(new_n915), .C2(new_n623), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n915), .B2(new_n640), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n354), .A3(new_n661), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


