//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  NOR3_X1   g046(.A1(new_n463), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT68), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(new_n478), .B2(new_n462), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n480));
  INV_X1    g055(.A(G100), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(new_n462), .ZN(new_n482));
  INV_X1    g057(.A(new_n476), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n462), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n482), .B(new_n487), .C1(G124), .C2(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n465), .A3(G2104), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n475), .A2(new_n492), .A3(G126), .A4(new_n464), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT70), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(KEYINPUT70), .B2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n463), .A2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G102), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n464), .A2(new_n466), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR4_X1   g078(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n503), .A2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n475), .A2(new_n492), .A3(new_n464), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n475), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n500), .B1(new_n513), .B2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT74), .Z(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n519), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n522), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n530), .B(new_n532), .C1(new_n536), .C2(KEYINPUT75), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(KEYINPUT75), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  INV_X1    g114(.A(new_n523), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(G52), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n519), .A2(G64), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n516), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n540), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n531), .A2(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n550), .B(new_n551), .C1(new_n516), .C2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT77), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  AOI22_X1  g134(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n516), .B1(new_n523), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n531), .A2(G53), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n563), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n540), .A2(G87), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT79), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n519), .A2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(G651), .A2(new_n575), .B1(new_n531), .B2(G49), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G288));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n523), .A2(new_n578), .B1(new_n525), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n519), .A2(G61), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(KEYINPUT80), .B1(G73), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n519), .A2(new_n584), .A3(G61), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n516), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT81), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n588));
  AOI211_X1 g163(.A(new_n588), .B(new_n516), .C1(new_n583), .C2(new_n585), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n581), .B1(new_n587), .B2(new_n589), .ZN(G305));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n523), .A2(new_n591), .B1(new_n525), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n516), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n540), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(new_n519), .A2(G66), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n516), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G54), .B2(new_n531), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  XOR2_X1   g187(.A(KEYINPUT82), .B(G559), .Z(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(G860), .B2(new_n613), .ZN(G148));
  INV_X1    g189(.A(new_n554), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n606), .A2(G868), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT11), .Z(G282));
  INV_X1    g194(.A(new_n618), .ZN(G323));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n623));
  OAI22_X1  g198(.A1(new_n488), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G135), .B2(new_n485), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n467), .A2(new_n498), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  MUX2_X1   g231(.A(new_n653), .B(new_n648), .S(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n666), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n669));
  OAI221_X1 g244(.A(new_n665), .B1(new_n667), .B2(new_n661), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G24), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n596), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n672), .ZN(new_n682));
  NOR2_X1   g257(.A1(G25), .A2(G29), .ZN(new_n683));
  INV_X1    g258(.A(G119), .ZN(new_n684));
  NOR2_X1   g259(.A1(G95), .A2(G2105), .ZN(new_n685));
  OAI21_X1  g260(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n686));
  OAI22_X1  g261(.A1(new_n488), .A2(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G131), .B2(new_n485), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n683), .B1(new_n688), .B2(G29), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT35), .B(G1991), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n682), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n689), .B2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(G305), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G6), .B2(G16), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n679), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n679), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT33), .B(G1976), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n679), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n679), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n693), .B1(new_n710), .B2(KEYINPUT34), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT86), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT36), .Z(new_n715));
  INV_X1    g290(.A(KEYINPUT24), .ZN(new_n716));
  INV_X1    g291(.A(G34), .ZN(new_n717));
  AOI21_X1  g292(.A(G29), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(G160), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2084), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(G32), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT26), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n726), .A2(new_n727), .B1(G105), .B2(new_n498), .ZN(new_n728));
  INV_X1    g303(.A(G129), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n488), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G141), .B2(new_n485), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n723), .B1(new_n731), .B2(new_n720), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT27), .B(G1996), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n720), .A2(G33), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  INV_X1    g311(.A(G139), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n484), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(G115), .A2(G2104), .ZN(new_n742));
  INV_X1    g317(.A(G127), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n501), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n740), .A2(new_n741), .B1(G2105), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n734), .B1(new_n745), .B2(new_n720), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n722), .B1(new_n732), .B2(new_n733), .C1(new_n746), .C2(G2072), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G2072), .B2(new_n746), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT89), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n720), .A2(G35), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n720), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT29), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(G2090), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n720), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  INV_X1    g332(.A(G128), .ZN(new_n758));
  NOR2_X1   g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n488), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G140), .B2(new_n485), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(new_n720), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT87), .B(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n679), .A2(G19), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n554), .B2(new_n679), .ZN(new_n768));
  INV_X1    g343(.A(G1341), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n679), .A2(G4), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n606), .B2(new_n679), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G1348), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n625), .A2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT31), .B(G11), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n776), .A2(G28), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n720), .B1(new_n776), .B2(G28), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n774), .B(new_n775), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n772), .B2(G1348), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n766), .A2(new_n770), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n754), .A2(new_n755), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G171), .A2(new_n679), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G5), .B2(new_n679), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT91), .Z(new_n788));
  AOI22_X1  g363(.A1(new_n785), .A2(new_n786), .B1(new_n732), .B2(new_n733), .ZN(new_n789));
  NAND2_X1  g364(.A1(G286), .A2(G16), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n679), .A2(G21), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1966), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n793), .C1(G2084), .C2(new_n721), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(G1966), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT90), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n679), .A2(G20), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT23), .Z(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G299), .B2(G16), .ZN(new_n800));
  INV_X1    g375(.A(G1956), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G2078), .ZN(new_n805));
  NAND2_X1  g380(.A1(G164), .A2(G29), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G27), .B2(G29), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n805), .B2(new_n807), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n715), .A2(new_n749), .A3(new_n783), .A4(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  NAND2_X1  g386(.A1(new_n531), .A2(G55), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT93), .B(G93), .Z(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n516), .B2(new_n813), .C1(new_n523), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT94), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(new_n553), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n554), .A2(new_n815), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n817), .A2(KEYINPUT95), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT95), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT96), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n606), .A2(G559), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n823), .B(new_n824), .Z(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  INV_X1    g403(.A(new_n816), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n831), .ZN(G145));
  NAND2_X1  g407(.A1(new_n511), .A2(new_n512), .ZN(new_n833));
  INV_X1    g408(.A(new_n504), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n514), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n500), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n762), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n745), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(G106), .A2(G2105), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n488), .A2(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G142), .B2(new_n485), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n628), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n841), .B(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n625), .B(G160), .Z(new_n849));
  XNOR2_X1  g424(.A(G162), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n688), .B(new_n731), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT98), .B(G37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g432(.A1(new_n606), .A2(new_n613), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n821), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n606), .B(G299), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G299), .B(new_n605), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT41), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n859), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n859), .B2(new_n860), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  XNOR2_X1  g444(.A(G305), .B(G303), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(G288), .B(G290), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(KEYINPUT99), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(KEYINPUT99), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n874), .B2(new_n871), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n868), .A2(new_n869), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n868), .B2(new_n869), .ZN(new_n878));
  OAI21_X1  g453(.A(G868), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(G868), .B2(new_n816), .ZN(G295));
  OAI21_X1  g455(.A(new_n879), .B1(G868), .B2(new_n816), .ZN(G331));
  NAND2_X1  g456(.A1(new_n862), .A2(new_n864), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n819), .A2(new_n820), .A3(G171), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(G171), .B1(new_n819), .B2(new_n820), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(G168), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(G168), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n860), .A3(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n875), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n891), .A3(new_n876), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n854), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT100), .B1(new_n860), .B2(new_n861), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(new_n864), .Z(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n887), .B2(new_n888), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n876), .B1(new_n900), .B2(new_n891), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n903));
  MUX2_X1   g478(.A(new_n896), .B(new_n902), .S(new_n903), .Z(new_n904));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n897), .B2(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n900), .A2(new_n891), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n875), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(KEYINPUT101), .A3(new_n854), .A4(new_n895), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT43), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n893), .A2(new_n903), .A3(new_n894), .A4(new_n895), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n913), .A2(KEYINPUT44), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT102), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT102), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n906), .B1(new_n915), .B2(new_n916), .ZN(G397));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n837), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(G160), .A2(G40), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(G1996), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n731), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT104), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n923), .B(KEYINPUT105), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n762), .B(G2067), .ZN(new_n928));
  INV_X1    g503(.A(G1996), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n731), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n688), .A2(new_n690), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n688), .A2(new_n690), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n923), .A2(G1986), .A3(G290), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n923), .A2(new_n672), .A3(new_n596), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT103), .Z(new_n939));
  NOR2_X1   g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT106), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT107), .B1(G164), .B2(G1384), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n510), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT72), .B1(new_n509), .B2(new_n510), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(new_n504), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n943), .B(new_n918), .C1(new_n946), .C2(new_n500), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n942), .A2(new_n947), .A3(KEYINPUT108), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n921), .A2(G2090), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n837), .A2(KEYINPUT45), .A3(new_n918), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n920), .B1(G164), .B2(G1384), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(new_n922), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n955), .A2(new_n956), .B1(G1971), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n955), .A2(new_n956), .ZN(new_n961));
  OAI21_X1  g536(.A(G8), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G303), .A2(G8), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT55), .Z(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G305), .A2(G1981), .ZN(new_n967));
  INV_X1    g542(.A(G1981), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT110), .B1(new_n694), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  NOR3_X1   g545(.A1(G305), .A2(new_n970), .A3(G1981), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n942), .A2(new_n947), .A3(new_n922), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(G8), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT49), .B(new_n967), .C1(new_n969), .C2(new_n971), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n701), .A2(G1976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n975), .A2(G8), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT52), .ZN(new_n981));
  INV_X1    g556(.A(G1976), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n976), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT63), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(G8), .B(new_n964), .C1(new_n960), .C2(new_n961), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n966), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1966), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n942), .B2(new_n947), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n957), .A2(new_n922), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT112), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n921), .A2(G2084), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(G8), .A3(G168), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT113), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n990), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n978), .A2(new_n982), .A3(new_n701), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n969), .A2(new_n971), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n976), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n988), .B2(new_n985), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(KEYINPUT111), .C1(new_n988), .C2(new_n985), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1004), .A2(KEYINPUT63), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n948), .B1(new_n942), .B2(new_n947), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n922), .B1(new_n919), .B2(KEYINPUT50), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(G2090), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n959), .A2(G1971), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n985), .B1(new_n965), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n943), .B1(new_n837), .B2(new_n918), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT107), .B(G1384), .C1(new_n835), .C2(new_n836), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n920), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(G164), .A2(G1384), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n921), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n805), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(KEYINPUT118), .A3(new_n805), .A4(new_n1023), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(KEYINPUT53), .A3(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n957), .A2(new_n958), .A3(new_n805), .A4(new_n922), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n922), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT119), .B(G1961), .Z(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G301), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1018), .A2(new_n988), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n996), .B1(new_n1038), .B2(new_n991), .ZN(new_n1039));
  INV_X1    g614(.A(new_n997), .ZN(new_n1040));
  OAI211_X1 g615(.A(G168), .B(new_n1000), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(KEYINPUT117), .A3(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT51), .ZN(new_n1043));
  AOI21_X1  g618(.A(G168), .B1(new_n998), .B2(new_n1000), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  OAI211_X1 g621(.A(G8), .B(new_n1041), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1037), .B1(new_n1048), .B2(KEYINPUT62), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1049), .A2(KEYINPUT127), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT127), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1012), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1018), .A2(new_n988), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(KEYINPUT122), .B2(G2078), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n922), .B2(KEYINPUT121), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n921), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n957), .A2(new_n1062), .A3(new_n958), .A4(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1031), .A2(new_n1065), .A3(G301), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1058), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT123), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1057), .B1(new_n1071), .B2(new_n1036), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1028), .A2(new_n1035), .A3(G301), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1058), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1031), .A2(new_n1065), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT126), .B(G171), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(G301), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1057), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1056), .A2(new_n1072), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1348), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1033), .A2(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n975), .A2(G2067), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1085), .A3(KEYINPUT60), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n606), .A3(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1089), .A2(new_n606), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n562), .A2(KEYINPUT57), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n565), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT50), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n921), .B1(new_n1022), .B2(new_n948), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1956), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1023), .A2(new_n958), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1095), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT114), .B(new_n1095), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n801), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n959), .A2(new_n1099), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1094), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1103), .A2(KEYINPUT61), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT115), .B(G1996), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(new_n769), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n959), .A2(new_n1111), .B1(new_n975), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT59), .B1(new_n1114), .B2(new_n615), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n959), .A2(new_n1111), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n975), .A2(new_n1113), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1116), .B(new_n554), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1109), .A2(new_n1110), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1090), .A2(new_n1091), .A3(new_n1108), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1086), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n605), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1107), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1121), .A2(new_n1125), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1072), .A2(new_n1056), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1082), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1003), .B1(new_n966), .B2(new_n989), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1055), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n941), .B1(new_n1054), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n924), .B(KEYINPUT46), .Z(new_n1132));
  INV_X1    g707(.A(new_n927), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n928), .A2(new_n731), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT47), .Z(new_n1136));
  NAND2_X1  g711(.A1(new_n931), .A2(new_n932), .ZN(new_n1137));
  INV_X1    g712(.A(G2067), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n762), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1133), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n935), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n936), .B(KEYINPUT48), .Z(new_n1142));
  AOI211_X1 g717(.A(new_n1136), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1131), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g719(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n856), .A3(new_n1146), .ZN(G225));
  INV_X1    g721(.A(G225), .ZN(G308));
endmodule


