//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  INV_X1    g001(.A(G134gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G127gat), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT72), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n209), .A2(new_n217), .A3(KEYINPUT72), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n227), .C1(KEYINPUT69), .C2(KEYINPUT24), .ZN(new_n228));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  AND2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT69), .A2(KEYINPUT24), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n228), .A2(new_n230), .A3(new_n234), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n226), .A3(new_n227), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT24), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n232), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n246), .A2(new_n250), .A3(KEYINPUT66), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT66), .B1(new_n246), .B2(new_n250), .ZN(new_n252));
  AND4_X1   g051(.A1(KEYINPUT67), .A2(new_n237), .A3(new_n238), .A4(KEYINPUT23), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT67), .B1(new_n229), .B2(KEYINPUT23), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n240), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n256), .B2(KEYINPUT25), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n246), .A2(new_n250), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n246), .A2(new_n250), .A3(KEYINPUT66), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n230), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n229), .A2(KEYINPUT67), .A3(KEYINPUT23), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n263), .A2(new_n264), .B1(new_n239), .B2(new_n236), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n231), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n242), .B1(new_n257), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT27), .B(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n225), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n232), .B1(new_n270), .B2(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n239), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n229), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n277), .A3(new_n235), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n276), .B2(new_n229), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n273), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n223), .B1(new_n268), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n231), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT68), .B1(new_n266), .B2(new_n231), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n241), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n282), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n222), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G227gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT64), .Z(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G15gat), .B(G43gat), .Z(new_n297));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n292), .A2(KEYINPUT34), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n283), .B2(new_n288), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n283), .A2(new_n288), .ZN(new_n304));
  INV_X1    g103(.A(new_n291), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n303), .B1(new_n306), .B2(KEYINPUT34), .ZN(new_n307));
  INV_X1    g106(.A(new_n299), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n293), .B(KEYINPUT32), .C1(new_n295), .C2(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n300), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n300), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n202), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n300), .A2(new_n309), .ZN(new_n313));
  INV_X1    g112(.A(new_n307), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n307), .A3(new_n309), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(KEYINPUT81), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n321));
  INV_X1    g120(.A(G211gat), .ZN(new_n322));
  INV_X1    g121(.A(G218gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G226gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(new_n290), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n268), .A2(new_n282), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(KEYINPUT29), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n286), .B2(new_n287), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n331), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n268), .B2(new_n282), .ZN(new_n335));
  INV_X1    g134(.A(new_n329), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n286), .A2(new_n336), .A3(new_n287), .ZN(new_n337));
  INV_X1    g136(.A(new_n327), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND2_X1  g141(.A1(KEYINPUT73), .A2(KEYINPUT30), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(KEYINPUT73), .A2(KEYINPUT30), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n333), .A2(new_n339), .A3(new_n342), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n339), .ZN(new_n349));
  INV_X1    g148(.A(new_n342), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n339), .A3(new_n342), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  INV_X1    g156(.A(G155gat), .ZN(new_n358));
  INV_X1    g157(.A(G162gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G141gat), .B(G148gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n357), .B(new_n360), .C1(new_n361), .C2(KEYINPUT2), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G148gat), .ZN(new_n364));
  INV_X1    g163(.A(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G141gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n360), .A2(new_n357), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n357), .A2(KEYINPUT2), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n362), .A2(new_n209), .A3(new_n370), .A4(new_n217), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n362), .A2(new_n370), .B1(new_n209), .B2(new_n217), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n356), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n362), .A2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n218), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n371), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n356), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n354), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n362), .B2(new_n370), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n383), .A2(KEYINPUT74), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n362), .A2(new_n382), .A3(new_n370), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n385), .A2(new_n218), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(KEYINPUT74), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n376), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n220), .A2(new_n389), .A3(KEYINPUT4), .A4(new_n221), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n388), .A2(new_n355), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n385), .B(new_n218), .C1(new_n383), .C2(KEYINPUT74), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n383), .A2(KEYINPUT74), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n354), .B(new_n355), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n371), .A2(new_n391), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n220), .A2(new_n389), .A3(new_n221), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n391), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n381), .A2(new_n393), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402));
  XOR2_X1   g201(.A(G1gat), .B(G29gat), .Z(new_n403));
  XNOR2_X1  g202(.A(G57gat), .B(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n401), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n401), .A2(new_n410), .A3(new_n408), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n400), .A2(new_n388), .A3(new_n354), .A4(new_n355), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n379), .B1(new_n378), .B2(new_n356), .ZN(new_n413));
  AOI211_X1 g212(.A(KEYINPUT75), .B(new_n355), .C1(new_n377), .C2(new_n371), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT5), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n355), .B1(new_n394), .B2(new_n395), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n390), .A2(new_n392), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n412), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT78), .B1(new_n419), .B2(new_n407), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT6), .B1(new_n401), .B2(new_n408), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n409), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n319), .B1(new_n353), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G228gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n290), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n382), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n376), .ZN(new_n429));
  INV_X1    g228(.A(new_n385), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n327), .B1(new_n430), .B2(KEYINPUT29), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(G22gat), .A3(new_n431), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n427), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n434), .A2(new_n427), .A3(new_n435), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n440), .A2(KEYINPUT77), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n437), .B2(new_n443), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n335), .A2(new_n338), .A3(new_n337), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n338), .B1(new_n335), .B2(new_n337), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n350), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(new_n352), .A3(new_n344), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n410), .B1(new_n401), .B2(new_n408), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n419), .A2(KEYINPUT78), .A3(new_n407), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n422), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n409), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n456), .A2(new_n347), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n452), .B1(new_n461), .B2(KEYINPUT80), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n318), .A2(new_n424), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n315), .A2(new_n316), .A3(new_n450), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n456), .A2(new_n347), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n401), .A2(new_n408), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n402), .B1(new_n419), .B2(new_n407), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT35), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n450), .B1(new_n465), .B2(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(new_n449), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n444), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n355), .B1(new_n400), .B2(new_n388), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT39), .B1(new_n378), .B2(new_n356), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n407), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT40), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n420), .B(new_n411), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n473), .B1(new_n353), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n459), .A2(new_n460), .A3(new_n352), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n350), .B1(new_n349), .B2(KEYINPUT37), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n333), .B2(new_n339), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT38), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n350), .A2(KEYINPUT37), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n455), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n333), .A2(new_n492), .A3(new_n339), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT37), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n485), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n471), .B1(new_n484), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n310), .B2(new_n311), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n315), .A2(KEYINPUT36), .A3(new_n316), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n463), .A2(new_n470), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G197gat), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT11), .B(G169gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(G1gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT16), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G1gat), .B2(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G8gat), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n515), .B(new_n518), .C1(G1gat), .C2(new_n512), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G43gat), .ZN(new_n522));
  INV_X1    g321(.A(G50gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G43gat), .A2(G50gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n528));
  XOR2_X1   g327(.A(G43gat), .B(G50gat), .Z(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(KEYINPUT14), .ZN(new_n533));
  AND2_X1   g332(.A1(KEYINPUT83), .A2(G29gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(KEYINPUT83), .A2(G29gat), .ZN(new_n535));
  OAI21_X1  g334(.A(G36gat), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(KEYINPUT14), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n527), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(KEYINPUT84), .A2(KEYINPUT15), .ZN(new_n540));
  NOR2_X1   g339(.A1(KEYINPUT84), .A2(KEYINPUT15), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n524), .B(new_n525), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n527), .B1(new_n542), .B2(KEYINPUT85), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n521), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT13), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n539), .A2(new_n545), .A3(KEYINPUT17), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT17), .B1(new_n539), .B2(new_n545), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n521), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555));
  INV_X1    g354(.A(new_n546), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(new_n520), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n546), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n539), .A2(new_n545), .A3(KEYINPUT17), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n555), .A3(new_n521), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n551), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n550), .B1(new_n564), .B2(KEYINPUT18), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n566), .B(new_n551), .C1(new_n558), .C2(new_n563), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n511), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n558), .A2(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n548), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(KEYINPUT18), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n510), .A3(new_n572), .A4(new_n550), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT7), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n576), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(new_n585), .A3(new_n583), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n562), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT89), .Z(new_n592));
  INV_X1    g391(.A(KEYINPUT41), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n556), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n592), .A2(new_n593), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n203), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n359), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n597), .A2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n600), .A2(new_n605), .A3(new_n599), .A4(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G57gat), .B(G64gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT88), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n617), .A3(new_n611), .ZN(new_n618));
  INV_X1    g417(.A(new_n611), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT88), .B1(new_n619), .B2(new_n612), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n611), .A2(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G64gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(G57gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(KEYINPUT87), .A2(G57gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(KEYINPUT87), .A2(G57gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n628), .B2(G64gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n616), .B1(new_n622), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n520), .B1(new_n631), .B2(KEYINPUT21), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G231gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n290), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n631), .A2(KEYINPUT21), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(new_n631), .B2(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G127gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n205), .A3(new_n637), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n633), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n633), .A3(new_n640), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n358), .ZN(new_n645));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  AND3_X1   g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n610), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT92), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n589), .A2(new_n630), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT87), .B(G57gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n624), .B1(new_n654), .B2(new_n623), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n655), .A2(new_n618), .A3(new_n621), .A4(new_n620), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n656), .A2(new_n587), .A3(new_n588), .A4(new_n616), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n595), .A2(new_n631), .A3(KEYINPUT10), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n653), .B2(new_n657), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n652), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n674), .A2(new_n652), .A3(new_n666), .A4(new_n672), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n668), .A2(new_n672), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n651), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n504), .A2(new_n575), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n468), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  NOR4_X1   g484(.A1(new_n504), .A2(new_n465), .A3(new_n575), .A4(new_n681), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n518), .B2(new_n686), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT93), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n682), .A2(new_n695), .A3(new_n318), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT94), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n310), .A2(new_n311), .A3(new_n500), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT36), .B1(new_n315), .B2(new_n316), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT94), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n682), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n696), .B1(new_n703), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g503(.A1(new_n682), .A2(new_n473), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT95), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  OR2_X1    g507(.A1(new_n534), .A2(new_n535), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT98), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n711));
  NOR2_X1   g510(.A1(new_n609), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n700), .A2(new_n499), .A3(new_n701), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n310), .A2(new_n311), .A3(new_n473), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n353), .A2(new_n683), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n451), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n459), .A2(new_n460), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n465), .A2(KEYINPUT80), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n452), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n424), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n716), .B1(new_n720), .B2(new_n318), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n710), .B(new_n712), .C1(new_n713), .C2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n504), .B2(new_n609), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n463), .A2(new_n470), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n700), .A2(new_n499), .A3(new_n701), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n710), .B1(new_n727), .B2(new_n712), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n650), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n575), .A3(new_n679), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT96), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n709), .B1(new_n733), .B2(new_n468), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n504), .A2(new_n609), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(new_n731), .ZN(new_n736));
  INV_X1    g535(.A(new_n709), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n683), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(G1328gat));
  INV_X1    g539(.A(KEYINPUT99), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n733), .B2(new_n465), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n729), .A2(KEYINPUT99), .A3(new_n353), .A4(new_n732), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(G36gat), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(G36gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n736), .A2(new_n745), .A3(new_n353), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1329gat));
  OAI211_X1 g547(.A(new_n702), .B(new_n732), .C1(new_n724), .C2(new_n728), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G43gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n522), .A3(new_n318), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n749), .A2(G43gat), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n754), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n753), .A2(new_n755), .B1(KEYINPUT47), .B2(new_n757), .ZN(G1330gat));
  OAI211_X1 g557(.A(new_n473), .B(new_n732), .C1(new_n724), .C2(new_n728), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n450), .A2(G50gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT101), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n759), .A2(G50gat), .B1(new_n736), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT102), .A2(KEYINPUT48), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n762), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n768), .ZN(G1331gat));
  NOR4_X1   g568(.A1(new_n610), .A2(new_n650), .A3(new_n574), .A4(new_n680), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n727), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n468), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n628), .ZN(G1332gat));
  NOR2_X1   g572(.A1(new_n771), .A2(new_n465), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  INV_X1    g577(.A(new_n702), .ZN(new_n779));
  OAI21_X1  g578(.A(G71gat), .B1(new_n771), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(G71gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n318), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n771), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g583(.A1(new_n771), .A2(new_n450), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g585(.A1(new_n575), .A2(new_n650), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT103), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n680), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n729), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n576), .B1(new_n790), .B2(new_n683), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n788), .A2(new_n609), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT51), .B1(new_n727), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n792), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n680), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n796), .A2(new_n576), .A3(new_n683), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n791), .A2(new_n797), .ZN(G1336gat));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n577), .A3(new_n353), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n353), .B(new_n789), .C1(new_n724), .C2(new_n728), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G92gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g602(.A(G99gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(new_n804), .A3(new_n318), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n702), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n807), .B2(new_n804), .ZN(G1338gat));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n473), .B(new_n789), .C1(new_n724), .C2(new_n728), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n795), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n450), .A2(new_n680), .A3(G106gat), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT104), .Z(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n809), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n792), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n813), .B1(new_n817), .B2(new_n793), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n809), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(G106gat), .B2(new_n810), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT105), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n812), .B2(new_n813), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT105), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n810), .A2(G106gat), .B1(new_n812), .B2(new_n814), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n809), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(KEYINPUT106), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n659), .A2(new_n660), .A3(new_n663), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n671), .B1(new_n674), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n674), .A2(new_n666), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT92), .B1(new_n834), .B2(new_n671), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n835), .B2(new_n675), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT55), .B1(new_n830), .B2(new_n832), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n837), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n677), .A2(new_n839), .A3(KEYINPUT106), .A4(new_n833), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n574), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  OAI22_X1  g640(.A1(new_n569), .A2(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n508), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n679), .A2(new_n573), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n610), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n838), .A2(new_n840), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n573), .A2(new_n843), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n609), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n650), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n651), .A2(new_n575), .A3(new_n680), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT107), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT107), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NOR4_X1   g654(.A1(new_n855), .A2(new_n468), .A3(new_n353), .A4(new_n464), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT108), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n212), .A3(new_n574), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n855), .A2(new_n473), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(new_n683), .A3(new_n465), .A4(new_n318), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n575), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n210), .A3(new_n679), .ZN(new_n863));
  OAI21_X1  g662(.A(G120gat), .B1(new_n860), .B2(new_n680), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n860), .B2(new_n650), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n856), .A2(new_n205), .A3(new_n730), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT109), .ZN(G1342gat));
  NAND3_X1  g668(.A1(new_n856), .A2(new_n203), .A3(new_n610), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n860), .B2(new_n609), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n852), .A2(new_n875), .A3(new_n473), .A4(new_n854), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n702), .A2(new_n468), .A3(new_n353), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT110), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n844), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n830), .A2(new_n832), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n836), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n574), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n679), .A2(new_n573), .A3(new_n843), .A4(KEYINPUT110), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n609), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n848), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n879), .A2(new_n844), .B1(new_n883), .B2(new_n574), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n610), .B1(new_n890), .B2(new_n885), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT113), .A3(new_n650), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n850), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n730), .B1(new_n889), .B2(new_n892), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(KEYINPUT113), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n473), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n878), .B1(new_n898), .B2(KEYINPUT57), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n363), .B1(new_n899), .B2(new_n574), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n779), .A2(new_n473), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n855), .A2(new_n901), .A3(new_n468), .A4(new_n353), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n363), .A3(new_n574), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT58), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n878), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n896), .A2(KEYINPUT113), .ZN(new_n907));
  INV_X1    g706(.A(new_n850), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n896), .B2(KEYINPUT113), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n450), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n906), .B1(new_n910), .B2(new_n875), .ZN(new_n911));
  OAI21_X1  g710(.A(G141gat), .B1(new_n911), .B2(new_n575), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n903), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n905), .A2(new_n914), .ZN(G1344gat));
  NOR2_X1   g714(.A1(new_n609), .A2(new_n847), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n836), .A2(new_n837), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n650), .B1(new_n891), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n450), .B1(new_n920), .B2(new_n850), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT115), .B1(new_n921), .B2(KEYINPUT57), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n887), .A2(new_n918), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n908), .B1(new_n924), .B2(new_n650), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n875), .C1(new_n925), .C2(new_n450), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n852), .A2(KEYINPUT57), .A3(new_n473), .A4(new_n854), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT114), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n679), .A3(new_n877), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n902), .A2(new_n365), .A3(new_n679), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n365), .B1(new_n899), .B2(new_n679), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(KEYINPUT59), .C2(new_n936), .ZN(G1345gat));
  AOI21_X1  g736(.A(G155gat), .B1(new_n902), .B2(new_n730), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n650), .A2(new_n358), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT116), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n899), .B2(new_n940), .ZN(G1346gat));
  AOI21_X1  g740(.A(G162gat), .B1(new_n902), .B2(new_n610), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n609), .A2(new_n359), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n899), .B2(new_n943), .ZN(G1347gat));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n855), .A2(new_n683), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n464), .A2(new_n465), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n575), .A2(G169gat), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n945), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n946), .A2(KEYINPUT117), .A3(new_n947), .A4(new_n949), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n683), .A2(new_n465), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n318), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT118), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n859), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957), .B2(new_n575), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(KEYINPUT119), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1348gat));
  OAI21_X1  g762(.A(new_n238), .B1(new_n948), .B2(new_n680), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT120), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n957), .A2(new_n238), .A3(new_n680), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n730), .A2(new_n269), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n948), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n969), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n946), .A2(KEYINPUT121), .A3(new_n947), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(G183gat), .B1(new_n957), .B2(new_n650), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT60), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT60), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n973), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1350gat));
  NAND4_X1  g778(.A1(new_n946), .A2(new_n225), .A3(new_n610), .A4(new_n947), .ZN(new_n980));
  OAI21_X1  g779(.A(G190gat), .B1(new_n957), .B2(new_n609), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT122), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n984), .B(G190gat), .C1(new_n957), .C2(new_n609), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n983), .B1(new_n982), .B2(new_n985), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(G1351gat));
  NOR2_X1   g787(.A1(new_n901), .A2(new_n465), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n946), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g789(.A(KEYINPUT123), .B(G197gat), .ZN(new_n991));
  OR3_X1    g790(.A1(new_n990), .A2(new_n575), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n779), .A2(new_n954), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n849), .A2(new_n853), .A3(new_n850), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n853), .B1(new_n849), .B2(new_n850), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n996), .A2(KEYINPUT114), .A3(KEYINPUT57), .A4(new_n473), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n928), .A2(new_n929), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n993), .B1(new_n999), .B2(new_n927), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(new_n1001), .A3(new_n574), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(new_n991), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1001), .B1(new_n1000), .B2(new_n574), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n992), .B1(new_n1003), .B2(new_n1004), .ZN(G1352gat));
  NOR3_X1   g804(.A1(new_n990), .A2(G204gat), .A3(new_n680), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1006), .B1(KEYINPUT125), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g807(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1000), .A2(new_n679), .ZN(new_n1010));
  INV_X1    g809(.A(G204gat), .ZN(new_n1011));
  OAI221_X1 g810(.A(new_n1008), .B1(new_n1006), .B2(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(G1353gat));
  NAND4_X1  g811(.A1(new_n946), .A2(new_n322), .A3(new_n730), .A4(new_n989), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT63), .ZN(new_n1014));
  AOI211_X1 g813(.A(new_n1014), .B(new_n322), .C1(new_n1000), .C2(new_n730), .ZN(new_n1015));
  INV_X1    g814(.A(new_n993), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n932), .A2(new_n730), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(KEYINPUT63), .B1(new_n1017), .B2(G211gat), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1013), .B1(new_n1015), .B2(new_n1018), .ZN(G1354gat));
  NAND3_X1  g818(.A1(new_n946), .A2(new_n610), .A3(new_n989), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(new_n323), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1022));
  XNOR2_X1  g821(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1024));
  AOI211_X1 g823(.A(new_n323), .B(new_n609), .C1(new_n1000), .C2(new_n1024), .ZN(new_n1025));
  OR2_X1    g824(.A1(new_n1000), .A2(new_n1024), .ZN(new_n1026));
  AOI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1355gat));
endmodule


