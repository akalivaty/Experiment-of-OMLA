

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U558 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U559 ( .A1(n716), .A2(n983), .ZN(n709) );
  NOR2_X1 U560 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U561 ( .A(n729), .B(n728), .ZN(n735) );
  INV_X1 U562 ( .A(KEYINPUT102), .ZN(n708) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n728) );
  NOR2_X1 U564 ( .A1(G2084), .A2(n747), .ZN(n736) );
  INV_X1 U565 ( .A(KEYINPUT12), .ZN(n581) );
  XNOR2_X1 U566 ( .A(n581), .B(KEYINPUT71), .ZN(n582) );
  XNOR2_X1 U567 ( .A(n583), .B(n582), .ZN(n585) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n805) );
  NOR2_X1 U569 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  NOR2_X1 U571 ( .A1(n820), .A2(n819), .ZN(n822) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n652) );
  NOR2_X1 U573 ( .A1(G651), .A2(n642), .ZN(n662) );
  XOR2_X1 U574 ( .A(KEYINPUT17), .B(n525), .Z(n888) );
  NAND2_X1 U575 ( .A1(n888), .A2(G138), .ZN(n527) );
  INV_X1 U576 ( .A(G2105), .ZN(n528) );
  AND2_X1 U577 ( .A1(n528), .A2(G2104), .ZN(n889) );
  NAND2_X1 U578 ( .A1(G102), .A2(n889), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n532) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NAND2_X1 U581 ( .A1(G114), .A2(n894), .ZN(n530) );
  NOR2_X1 U582 ( .A1(G2104), .A2(n528), .ZN(n892) );
  NAND2_X1 U583 ( .A1(G126), .A2(n892), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(G164) );
  XOR2_X1 U586 ( .A(G2438), .B(G2454), .Z(n534) );
  XNOR2_X1 U587 ( .A(G2435), .B(G2430), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U589 ( .A(n535), .B(G2427), .Z(n537) );
  XNOR2_X1 U590 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U591 ( .A(n537), .B(n536), .ZN(n541) );
  XOR2_X1 U592 ( .A(G2443), .B(G2446), .Z(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT108), .B(G2451), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U595 ( .A(n541), .B(n540), .Z(n542) );
  AND2_X1 U596 ( .A1(G14), .A2(n542), .ZN(G401) );
  XOR2_X1 U597 ( .A(KEYINPUT64), .B(G651), .Z(n548) );
  NOR2_X1 U598 ( .A1(G543), .A2(n548), .ZN(n543) );
  XOR2_X2 U599 ( .A(KEYINPUT1), .B(n543), .Z(n653) );
  NAND2_X1 U600 ( .A1(n653), .A2(G64), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT66), .ZN(n547) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  NAND2_X1 U603 ( .A1(G52), .A2(n662), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT67), .B(n545), .Z(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G90), .A2(n652), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n642), .A2(n548), .ZN(n657) );
  NAND2_X1 U608 ( .A1(G77), .A2(n657), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U611 ( .A1(n553), .A2(n552), .ZN(G171) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U613 ( .A1(G135), .A2(n888), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G111), .A2(n894), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n892), .A2(G123), .ZN(n556) );
  XOR2_X1 U617 ( .A(KEYINPUT18), .B(n556), .Z(n557) );
  NOR2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n889), .A2(G99), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n934) );
  XNOR2_X1 U621 ( .A(G2096), .B(n934), .ZN(n561) );
  OR2_X1 U622 ( .A1(G2100), .A2(n561), .ZN(G156) );
  INV_X1 U623 ( .A(G108), .ZN(G238) );
  INV_X1 U624 ( .A(G120), .ZN(G236) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  NAND2_X1 U626 ( .A1(G63), .A2(n653), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT79), .B(n562), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n662), .A2(G51), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT80), .B(n563), .Z(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT6), .B(n566), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G76), .A2(n657), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT77), .B(n567), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n652), .A2(G89), .ZN(n568) );
  XOR2_X1 U635 ( .A(n568), .B(KEYINPUT4), .Z(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT5), .B(n571), .Z(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT78), .B(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT7), .B(n575), .ZN(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U642 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n577) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(G223) );
  INV_X1 U645 ( .A(G567), .ZN(n691) );
  NOR2_X1 U646 ( .A1(n691), .A2(G223), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n578), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U648 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n580) );
  NAND2_X1 U649 ( .A1(G56), .A2(n653), .ZN(n579) );
  XNOR2_X1 U650 ( .A(n580), .B(n579), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G81), .A2(n652), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G68), .A2(n657), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U654 ( .A(KEYINPUT13), .B(n586), .Z(n587) );
  XNOR2_X1 U655 ( .A(n589), .B(KEYINPUT72), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G43), .A2(n662), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n987) );
  INV_X1 U658 ( .A(G860), .ZN(n614) );
  OR2_X1 U659 ( .A1(n987), .A2(n614), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT73), .B(n592), .Z(G153) );
  INV_X1 U661 ( .A(G171), .ZN(G301) );
  NAND2_X1 U662 ( .A1(n652), .A2(G92), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G66), .A2(n653), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n662), .A2(G54), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G79), .A2(n657), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U668 ( .A(KEYINPUT75), .B(n597), .Z(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U670 ( .A(KEYINPUT15), .B(n600), .ZN(n983) );
  INV_X1 U671 ( .A(G868), .ZN(n673) );
  NAND2_X1 U672 ( .A1(n983), .A2(n673), .ZN(n601) );
  XNOR2_X1 U673 ( .A(KEYINPUT76), .B(n601), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G868), .A2(G301), .ZN(n602) );
  XNOR2_X1 U675 ( .A(KEYINPUT74), .B(n602), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U677 ( .A1(G91), .A2(n652), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G53), .A2(n662), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n657), .A2(G78), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT68), .B(n607), .Z(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G65), .A2(n653), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G299) );
  NOR2_X1 U685 ( .A1(G286), .A2(n673), .ZN(n613) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n614), .A2(G559), .ZN(n615) );
  INV_X1 U689 ( .A(n983), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n615), .A2(n621), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(n983), .A2(n673), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT81), .ZN(n618) );
  NOR2_X1 U694 ( .A1(G559), .A2(n618), .ZN(n620) );
  NOR2_X1 U695 ( .A1(G868), .A2(n987), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U697 ( .A1(n621), .A2(G559), .ZN(n671) );
  XNOR2_X1 U698 ( .A(n987), .B(n671), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n622), .A2(G860), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G93), .A2(n652), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT82), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G67), .A2(n653), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n662), .A2(G55), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G80), .A2(n657), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n674) );
  XOR2_X1 U708 ( .A(n630), .B(n674), .Z(G145) );
  NAND2_X1 U709 ( .A1(G62), .A2(n653), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G75), .A2(n657), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n652), .A2(G88), .ZN(n633) );
  XOR2_X1 U713 ( .A(KEYINPUT86), .B(n633), .Z(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n662), .A2(G50), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(G303) );
  NAND2_X1 U717 ( .A1(G49), .A2(n662), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n653), .A2(n640), .ZN(n641) );
  XOR2_X1 U721 ( .A(KEYINPUT83), .B(n641), .Z(n644) );
  NAND2_X1 U722 ( .A1(n642), .A2(G87), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U724 ( .A1(n662), .A2(G47), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G60), .A2(n653), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U727 ( .A(KEYINPUT65), .B(n647), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n657), .A2(G72), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G85), .A2(n652), .ZN(n648) );
  AND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(G290) );
  NAND2_X1 U732 ( .A1(n652), .A2(G86), .ZN(n655) );
  NAND2_X1 U733 ( .A1(G61), .A2(n653), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U735 ( .A(KEYINPUT84), .B(n656), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n657), .A2(G73), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(KEYINPUT2), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(KEYINPUT85), .ZN(n660) );
  NOR2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n662), .A2(G48), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(G305) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(G303), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n666), .B(G290), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(G305), .ZN(n668) );
  XOR2_X1 U746 ( .A(n674), .B(n668), .Z(n670) );
  INV_X1 U747 ( .A(G299), .ZN(n974) );
  XNOR2_X1 U748 ( .A(n987), .B(n974), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n911) );
  XOR2_X1 U750 ( .A(n911), .B(n671), .Z(n672) );
  NAND2_X1 U751 ( .A1(G868), .A2(n672), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n680), .A2(G2072), .ZN(n681) );
  XOR2_X1 U759 ( .A(KEYINPUT87), .B(n681), .Z(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U761 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n683) );
  NAND2_X1 U762 ( .A1(G132), .A2(G82), .ZN(n682) );
  XNOR2_X1 U763 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U764 ( .A(n684), .B(KEYINPUT88), .ZN(n685) );
  NOR2_X1 U765 ( .A1(G218), .A2(n685), .ZN(n686) );
  XNOR2_X1 U766 ( .A(KEYINPUT90), .B(n686), .ZN(n687) );
  NAND2_X1 U767 ( .A1(n687), .A2(G96), .ZN(n843) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n843), .ZN(n688) );
  XNOR2_X1 U769 ( .A(n688), .B(KEYINPUT91), .ZN(n693) );
  NOR2_X1 U770 ( .A1(G236), .A2(G238), .ZN(n689) );
  NAND2_X1 U771 ( .A1(G69), .A2(n689), .ZN(n690) );
  NOR2_X1 U772 ( .A1(G237), .A2(n690), .ZN(n845) );
  NOR2_X1 U773 ( .A1(n691), .A2(n845), .ZN(n692) );
  NOR2_X1 U774 ( .A1(n693), .A2(n692), .ZN(G319) );
  INV_X1 U775 ( .A(G319), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U777 ( .A1(n695), .A2(n694), .ZN(n842) );
  NAND2_X1 U778 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U779 ( .A1(n888), .A2(G137), .ZN(n698) );
  NAND2_X1 U780 ( .A1(G101), .A2(n889), .ZN(n696) );
  XOR2_X1 U781 ( .A(KEYINPUT23), .B(n696), .Z(n697) );
  NAND2_X1 U782 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U783 ( .A1(G113), .A2(n894), .ZN(n700) );
  NAND2_X1 U784 ( .A1(G125), .A2(n892), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U786 ( .A1(n702), .A2(n701), .ZN(G160) );
  INV_X1 U787 ( .A(G303), .ZN(G166) );
  NAND2_X1 U788 ( .A1(G160), .A2(G40), .ZN(n804) );
  INV_X1 U789 ( .A(n804), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n805), .A2(n703), .ZN(n747) );
  XNOR2_X1 U791 ( .A(G1996), .B(KEYINPUT101), .ZN(n949) );
  NOR2_X1 U792 ( .A1(n747), .A2(n949), .ZN(n704) );
  XNOR2_X1 U793 ( .A(n704), .B(KEYINPUT26), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n987), .A2(n705), .ZN(n707) );
  NAND2_X1 U795 ( .A1(G1341), .A2(n747), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n716) );
  XNOR2_X1 U797 ( .A(n709), .B(n708), .ZN(n715) );
  INV_X1 U798 ( .A(n747), .ZN(n730) );
  NAND2_X1 U799 ( .A1(G2067), .A2(n730), .ZN(n710) );
  XOR2_X1 U800 ( .A(KEYINPUT103), .B(n710), .Z(n712) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n747), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U803 ( .A(KEYINPUT104), .B(n713), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n716), .A2(n983), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n723) );
  NAND2_X1 U807 ( .A1(n730), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U808 ( .A(n719), .B(KEYINPUT27), .ZN(n721) );
  XOR2_X1 U809 ( .A(G1956), .B(KEYINPUT100), .Z(n998) );
  NOR2_X1 U810 ( .A1(n730), .A2(n998), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n974), .A2(n724), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U814 ( .A1(n974), .A2(n724), .ZN(n725) );
  XOR2_X1 U815 ( .A(n725), .B(KEYINPUT28), .Z(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n729) );
  OR2_X1 U817 ( .A1(n730), .A2(G1961), .ZN(n732) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U819 ( .A1(n730), .A2(n955), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n740) );
  AND2_X1 U821 ( .A1(n740), .A2(G171), .ZN(n733) );
  XNOR2_X1 U822 ( .A(n733), .B(KEYINPUT99), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n745) );
  NAND2_X1 U824 ( .A1(G8), .A2(n747), .ZN(n782) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n782), .ZN(n760) );
  XOR2_X1 U826 ( .A(KEYINPUT98), .B(n736), .Z(n756) );
  NAND2_X1 U827 ( .A1(G8), .A2(n756), .ZN(n737) );
  NOR2_X1 U828 ( .A1(n760), .A2(n737), .ZN(n738) );
  XOR2_X1 U829 ( .A(KEYINPUT30), .B(n738), .Z(n739) );
  NOR2_X1 U830 ( .A1(G168), .A2(n739), .ZN(n742) );
  NOR2_X1 U831 ( .A1(G171), .A2(n740), .ZN(n741) );
  XOR2_X1 U832 ( .A(KEYINPUT31), .B(n743), .Z(n744) );
  NAND2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n758) );
  NAND2_X1 U834 ( .A1(n758), .A2(G286), .ZN(n754) );
  INV_X1 U835 ( .A(G8), .ZN(n752) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n782), .ZN(n746) );
  XNOR2_X1 U837 ( .A(KEYINPUT105), .B(n746), .ZN(n750) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U839 ( .A1(G166), .A2(n748), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  OR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U843 ( .A(n755), .B(KEYINPUT32), .ZN(n764) );
  INV_X1 U844 ( .A(n756), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n757), .A2(G8), .ZN(n762) );
  INV_X1 U846 ( .A(n758), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n764), .A2(n763), .ZN(n778) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n771) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n771), .A2(n765), .ZN(n975) );
  NAND2_X1 U853 ( .A1(n778), .A2(n975), .ZN(n768) );
  INV_X1 U854 ( .A(n782), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n973) );
  AND2_X1 U856 ( .A1(n766), .A2(n973), .ZN(n767) );
  AND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U858 ( .A1(n769), .A2(KEYINPUT33), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT106), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n771), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n782), .A2(n772), .ZN(n773) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n969) );
  NAND2_X1 U863 ( .A1(n775), .A2(n969), .ZN(n786) );
  NOR2_X1 U864 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n779), .A2(n782), .ZN(n784) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U869 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  OR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  AND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n820) );
  NAND2_X1 U873 ( .A1(G141), .A2(n888), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G117), .A2(n894), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n889), .A2(G105), .ZN(n789) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n789), .Z(n790) );
  NOR2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n892), .A2(G129), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n903) );
  NAND2_X1 U881 ( .A1(G1996), .A2(n903), .ZN(n803) );
  NAND2_X1 U882 ( .A1(G119), .A2(n892), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n794), .B(KEYINPUT94), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G95), .A2(n889), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G107), .A2(n894), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G131), .A2(n888), .ZN(n797) );
  XNOR2_X1 U888 ( .A(KEYINPUT95), .B(n797), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n876) );
  NAND2_X1 U891 ( .A1(G1991), .A2(n876), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n925) );
  NOR2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n833) );
  NAND2_X1 U894 ( .A1(n925), .A2(n833), .ZN(n806) );
  XOR2_X1 U895 ( .A(KEYINPUT96), .B(n806), .Z(n825) );
  XNOR2_X1 U896 ( .A(KEYINPUT97), .B(n825), .ZN(n818) );
  NAND2_X1 U897 ( .A1(G116), .A2(n894), .ZN(n808) );
  NAND2_X1 U898 ( .A1(G128), .A2(n892), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U900 ( .A(KEYINPUT35), .B(n809), .Z(n816) );
  XNOR2_X1 U901 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n810) );
  XNOR2_X1 U902 ( .A(n810), .B(KEYINPUT34), .ZN(n814) );
  NAND2_X1 U903 ( .A1(G140), .A2(n888), .ZN(n812) );
  NAND2_X1 U904 ( .A1(G104), .A2(n889), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U906 ( .A(n814), .B(n813), .Z(n815) );
  NOR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n817), .ZN(n908) );
  XNOR2_X1 U909 ( .A(G2067), .B(KEYINPUT37), .ZN(n831) );
  NOR2_X1 U910 ( .A1(n908), .A2(n831), .ZN(n933) );
  NAND2_X1 U911 ( .A1(n833), .A2(n933), .ZN(n829) );
  NAND2_X1 U912 ( .A1(n818), .A2(n829), .ZN(n819) );
  XNOR2_X1 U913 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U914 ( .A1(n982), .A2(n833), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n836) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n903), .ZN(n930) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n876), .ZN(n936) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n936), .A2(n823), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n930), .A2(n826), .ZN(n828) );
  XOR2_X1 U922 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n908), .A2(n831), .ZN(n924) );
  NAND2_X1 U926 ( .A1(n832), .A2(n924), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n837), .ZN(G329) );
  INV_X1 U930 ( .A(G223), .ZN(n838) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U933 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  XOR2_X1 U935 ( .A(KEYINPUT109), .B(n840), .Z(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U938 ( .A(G132), .ZN(G219) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G82), .ZN(G220) );
  INV_X1 U941 ( .A(n843), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(G261) );
  INV_X1 U943 ( .A(G261), .ZN(G325) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2678), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT42), .B(G2090), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2096), .B(G2100), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U953 ( .A(G2078), .B(G2084), .Z(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1981), .B(G1966), .Z(n857) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n867) );
  XOR2_X1 U958 ( .A(G2474), .B(KEYINPUT41), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1961), .B(KEYINPUT114), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(G1976), .B(G1971), .Z(n861) );
  XNOR2_X1 U962 ( .A(G1986), .B(G1956), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G124), .A2(n892), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  XNOR2_X1 U970 ( .A(n869), .B(KEYINPUT115), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G112), .A2(n894), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G136), .A2(n888), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G100), .A2(n889), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT117), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U980 ( .A(G164), .B(n879), .ZN(n907) );
  NAND2_X1 U981 ( .A1(G118), .A2(n894), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G130), .A2(n892), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G142), .A2(n888), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G106), .A2(n889), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  XNOR2_X1 U988 ( .A(KEYINPUT116), .B(n885), .ZN(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n902) );
  NAND2_X1 U990 ( .A1(G139), .A2(n888), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n899) );
  NAND2_X1 U993 ( .A1(n892), .A2(G127), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n893), .B(KEYINPUT118), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n920) );
  XOR2_X1 U999 ( .A(G160), .B(n920), .Z(n900) );
  XNOR2_X1 U1000 ( .A(n934), .B(n900), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n903), .B(G162), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(G171), .B(G286), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(n913), .B(n983), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n916), .ZN(n917) );
  AND2_X1 U1014 ( .A1(G319), .A2(n917), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1019 ( .A(G2072), .B(n920), .Z(n922) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n923), .ZN(n928) );
  INV_X1 U1023 ( .A(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n942) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT51), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(G160), .B(G2084), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT119), .B(n938), .Z(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n943), .ZN(n944) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n965) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n965), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n960) );
  XNOR2_X1 U1041 ( .A(G1991), .B(G25), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n952) );
  XOR2_X1 U1046 ( .A(G32), .B(n949), .Z(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1050 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n967) );
  INV_X1 U1058 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n968), .ZN(n1024) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n993) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n971), .B(KEYINPUT57), .ZN(n991) );
  XNOR2_X1 U1065 ( .A(G171), .B(G1961), .ZN(n980) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n974), .B(G1956), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT121), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n984), .B(n983), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1341), .B(n987), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n1022) );
  INV_X1 U1080 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .Z(n994) );
  XNOR2_X1 U1082 ( .A(G4), .B(n994), .ZN(n1003) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1086 ( .A(KEYINPUT122), .B(n997), .Z(n1000) );
  XOR2_X1 U1087 ( .A(n998), .B(G20), .Z(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(n1001), .B(KEYINPUT123), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1004), .ZN(n1015) );
  XNOR2_X1 U1092 ( .A(G1966), .B(KEYINPUT124), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(n1005), .B(G21), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1986), .B(KEYINPUT125), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(G24), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  XOR2_X1 U1111 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

