//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT68), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT69), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n472), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n468), .A2(new_n469), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n468), .B2(new_n469), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(new_n490), .C1(new_n468), .C2(new_n469), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n461), .C1(new_n468), .C2(new_n469), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n464), .A2(new_n498), .A3(G138), .A4(new_n461), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT73), .A2(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT73), .A2(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g088(.A(KEYINPUT74), .B(G651), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT72), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n515), .A2(G88), .A3(new_n505), .A4(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n515), .A2(G50), .A3(G543), .A4(new_n517), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT75), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n508), .B1(new_n522), .B2(new_n523), .ZN(G166));
  AND3_X1   g099(.A1(new_n515), .A2(G543), .A3(new_n517), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n515), .A2(G89), .A3(new_n505), .A4(new_n517), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(new_n529), .A3(new_n532), .ZN(new_n534));
  NOR3_X1   g109(.A1(new_n528), .A2(new_n533), .A3(new_n534), .ZN(G168));
  NAND3_X1  g110(.A1(new_n515), .A2(new_n505), .A3(new_n517), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n525), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n507), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n525), .A2(G43), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n515), .A2(G81), .A3(new_n505), .A4(new_n517), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n507), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND4_X1  g129(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n517), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT78), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n525), .A2(new_n558), .A3(new_n559), .A4(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(new_n555), .B2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n555), .A2(new_n562), .A3(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n557), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n507), .B1(new_n565), .B2(KEYINPUT80), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n537), .A2(G91), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  AND3_X1   g145(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT75), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n518), .B2(new_n519), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n571), .A2(new_n572), .B1(new_n507), .B2(new_n506), .ZN(G303));
  NAND4_X1  g148(.A1(new_n515), .A2(G87), .A3(new_n505), .A4(new_n517), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G49), .A2(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n515), .A2(new_n517), .A3(new_n577), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND4_X1  g156(.A1(new_n515), .A2(G86), .A3(new_n505), .A4(new_n517), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n515), .A2(G48), .A3(G543), .A4(new_n517), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n505), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT82), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n525), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT83), .B(G85), .Z(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n507), .B2(new_n590), .C1(new_n536), .C2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n536), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n505), .A2(G66), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT84), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n525), .A2(G54), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT85), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  INV_X1    g188(.A(new_n548), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n608), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n604), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n464), .A2(new_n462), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT87), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n479), .A2(G135), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT88), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n481), .B2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  INV_X1    g208(.A(new_n632), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n622), .A2(new_n623), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n625), .A2(new_n633), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT89), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n623), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n635), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT90), .ZN(new_n670));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(KEYINPUT90), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n667), .A2(new_n668), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(new_n669), .ZN(new_n677));
  MUX2_X1   g252(.A(new_n677), .B(new_n676), .S(new_n672), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NOR2_X1   g261(.A1(G160), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(KEYINPUT24), .B2(G34), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(KEYINPUT24), .B2(G34), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G2084), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT99), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(G33), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n479), .A2(G139), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n464), .A2(G127), .ZN(new_n697));
  NAND2_X1  g272(.A1(G115), .A2(G2104), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n461), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT25), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n694), .B1(new_n702), .B2(new_n686), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G2072), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT101), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n479), .A2(G141), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n462), .A2(G105), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT26), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n709), .B(new_n711), .C1(G129), .C2(new_n481), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n686), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n686), .B2(G32), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n693), .B(new_n704), .C1(new_n706), .C2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G21), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G168), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT103), .B(G1966), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n717), .B(new_n718), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT105), .B(KEYINPUT23), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(G20), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G299), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1956), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT98), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n686), .A2(G26), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n481), .A2(G128), .ZN(new_n735));
  INV_X1    g310(.A(G140), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n465), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n738));
  INV_X1    g313(.A(G116), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n686), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G2067), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n715), .A2(new_n706), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n634), .A2(G29), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(KEYINPUT104), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G11), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT30), .B(G28), .Z(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n747), .B2(KEYINPUT104), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n745), .A2(new_n746), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n686), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n686), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G2090), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n687), .A2(G2084), .A3(new_n689), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n686), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n686), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n756), .B2(G2090), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n753), .A2(new_n757), .A3(new_n758), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G19), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n548), .B2(G16), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G1341), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(G1341), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n719), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n719), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(G1961), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n767), .B(new_n771), .C1(G1961), .C2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n719), .A2(G4), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n605), .B2(new_n719), .ZN(new_n774));
  INV_X1    g349(.A(G1348), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n721), .A2(new_n723), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n764), .A2(new_n772), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n724), .A2(new_n730), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(KEYINPUT94), .ZN(new_n782));
  OR2_X1    g357(.A1(G16), .A2(G23), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G288), .B2(new_n719), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT92), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(G6), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G305), .B2(new_n719), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n790), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n788), .B(new_n792), .C1(G305), .C2(new_n719), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n786), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(new_n783), .C1(G288), .C2(new_n719), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n787), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n719), .A2(G22), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G303), .B2(G16), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G1971), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G1971), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n797), .B(new_n798), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G290), .A2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G24), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(G16), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G1986), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n805), .B(G1986), .C1(G16), .C2(new_n806), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n479), .A2(G131), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n481), .A2(G119), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G29), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n818));
  OR2_X1    g393(.A1(G25), .A2(G29), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OR3_X1    g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n809), .A2(new_n810), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n804), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT93), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n804), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n787), .A2(new_n794), .A3(new_n796), .ZN(new_n831));
  INV_X1    g406(.A(new_n801), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n802), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n798), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n828), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n836), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n836), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n782), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n804), .A2(new_n829), .A3(new_n826), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n829), .B1(new_n804), .B2(new_n826), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n844), .A2(new_n845), .A3(new_n834), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT95), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  INV_X1    g422(.A(new_n782), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n836), .A2(new_n837), .A3(new_n840), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n780), .B1(new_n843), .B2(new_n850), .ZN(G311));
  NOR3_X1   g426(.A1(new_n841), .A2(new_n842), .A3(new_n782), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n779), .B1(new_n852), .B2(new_n853), .ZN(G150));
  NAND4_X1  g429(.A1(new_n515), .A2(G93), .A3(new_n505), .A4(new_n517), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n515), .A2(G55), .A3(G543), .A4(new_n517), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n855), .B(new_n856), .C1(new_n507), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n604), .A2(new_n612), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n858), .B(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n614), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n548), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n864), .B(new_n870), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  INV_X1    g447(.A(G860), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n871), .B2(KEYINPUT39), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n861), .B1(new_n872), .B2(new_n874), .ZN(G145));
  XNOR2_X1  g450(.A(G160), .B(new_n485), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n634), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n708), .A2(new_n712), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n501), .ZN(new_n881));
  INV_X1    g456(.A(new_n742), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n880), .A2(new_n501), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n501), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n742), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n481), .A2(G130), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT110), .Z(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(G118), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(G2105), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n479), .B2(G142), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n815), .B(new_n621), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n877), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(KEYINPUT111), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n883), .A2(new_n903), .A3(new_n886), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n883), .A2(new_n886), .A3(new_n903), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n883), .B2(new_n886), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n877), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT112), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n899), .B2(new_n904), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(KEYINPUT112), .A3(new_n908), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  NAND2_X1  g492(.A1(new_n858), .A2(new_n608), .ZN(new_n918));
  XNOR2_X1  g493(.A(G166), .B(G290), .ZN(new_n919));
  XNOR2_X1  g494(.A(G288), .B(G305), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT113), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(KEYINPUT113), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n870), .B(new_n616), .ZN(new_n925));
  NOR2_X1   g500(.A1(G299), .A2(new_n604), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G299), .A2(new_n604), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n924), .B(new_n930), .C1(new_n935), .C2(new_n925), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n935), .B2(new_n925), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(KEYINPUT113), .A3(new_n922), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n923), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n918), .B1(new_n939), .B2(new_n608), .ZN(G295));
  OAI21_X1  g515(.A(new_n918), .B1(new_n939), .B2(new_n608), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n867), .A2(new_n548), .A3(new_n868), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n548), .B1(new_n867), .B2(new_n868), .ZN(new_n944));
  OAI21_X1  g519(.A(G171), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n866), .A2(G301), .A3(new_n869), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G286), .ZN(new_n948));
  INV_X1    g523(.A(new_n929), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n946), .A3(G168), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n945), .A2(new_n946), .A3(G168), .ZN(new_n952));
  AOI21_X1  g527(.A(G168), .B1(new_n945), .B2(new_n946), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(new_n934), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n955), .B2(new_n921), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(new_n921), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n951), .B(new_n958), .C1(new_n954), .C2(new_n934), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n956), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n942), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n955), .A2(new_n921), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n909), .A3(new_n959), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT44), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(KEYINPUT120), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n501), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT50), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n495), .B2(new_n500), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT115), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(KEYINPUT114), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n976), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2090), .ZN(new_n983));
  INV_X1    g558(.A(new_n467), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT70), .B1(new_n472), .B2(G2105), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n474), .B(new_n461), .C1(new_n470), .C2(new_n471), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n984), .B(G40), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n978), .A2(new_n982), .A3(new_n983), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n972), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n975), .A2(KEYINPUT45), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1971), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n970), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G166), .B2(new_n970), .ZN(new_n998));
  NAND3_X1  g573(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT114), .B1(new_n501), .B2(new_n971), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n979), .B(G1384), .C1(new_n495), .C2(new_n500), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n988), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n576), .A2(new_n579), .A3(G1976), .A4(new_n580), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(G288), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n970), .B1(new_n1005), .B2(new_n988), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n1007), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G305), .A2(G1981), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n582), .A2(new_n583), .A3(new_n1015), .A4(new_n587), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT117), .B(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1012), .B(new_n1017), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1020), .A2(new_n1018), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1009), .B(new_n1013), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G288), .A2(G1976), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1016), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1002), .A2(new_n1024), .B1(new_n1027), .B2(new_n1012), .ZN(new_n1028));
  NOR3_X1   g603(.A1(G166), .A2(new_n997), .A3(new_n970), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n987), .B1(new_n976), .B2(new_n975), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n983), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n995), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(new_n1036), .A3(KEYINPUT119), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n970), .B1(new_n1034), .B2(new_n995), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1000), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT45), .B1(new_n980), .B2(new_n981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n988), .A2(new_n992), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n722), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n978), .A2(new_n982), .A3(new_n691), .A4(new_n988), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n970), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1046), .A2(G168), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1041), .A2(new_n1001), .A3(new_n1024), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT63), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1051));
  INV_X1    g626(.A(new_n996), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1031), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1002), .A2(new_n1023), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n969), .B(new_n1028), .C1(new_n1050), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT122), .B1(new_n1005), .B2(new_n988), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n1058));
  NOR4_X1   g633(.A1(new_n1003), .A2(new_n1004), .A3(new_n987), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n744), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n978), .A2(new_n982), .A3(new_n988), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n775), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n604), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1956), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n993), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n564), .A2(new_n568), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n564), .B2(new_n568), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1065), .B(new_n1069), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1063), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1070), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G299), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n564), .A2(new_n568), .A3(new_n1070), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1076), .B(new_n1077), .C1(new_n1064), .C2(new_n1068), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1073), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1060), .A2(new_n1062), .A3(new_n604), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1063), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1078), .A2(new_n1073), .A3(KEYINPUT61), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1006), .A2(new_n1058), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1005), .A2(KEYINPUT122), .A3(new_n988), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n993), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n614), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1060), .A2(new_n1062), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT123), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1096), .B(new_n1098), .C1(new_n1094), .C2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1079), .B1(new_n1086), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1044), .A2(new_n1045), .A3(G168), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G8), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(KEYINPUT124), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1104), .A2(new_n1106), .B1(G286), .B2(new_n1046), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(G8), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT53), .B1(new_n1091), .B2(new_n761), .ZN(new_n1111));
  INV_X1    g686(.A(G1961), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1061), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G301), .B(KEYINPUT54), .ZN(new_n1114));
  INV_X1    g689(.A(new_n992), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n975), .A2(KEYINPUT45), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT125), .B(G2078), .Z(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1119), .B(new_n467), .C1(G2105), .C2(new_n472), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1113), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1114), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1110), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1054), .A2(new_n1041), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1054), .A2(KEYINPUT126), .A3(new_n1041), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1102), .A2(new_n1127), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1048), .A2(new_n1049), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1028), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT120), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1046), .A2(G286), .ZN(new_n1138));
  AND4_X1   g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1109), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1125), .A2(G171), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1130), .A3(new_n1131), .A4(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1056), .A2(new_n1132), .A3(new_n1135), .A4(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n991), .A2(new_n987), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n742), .B(G2067), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n878), .B(new_n1092), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n816), .A2(new_n822), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n815), .A2(new_n823), .ZN(new_n1149));
  AND4_X1   g724(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G290), .A2(G1986), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(G290), .A2(G1986), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1145), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1144), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1145), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1147), .A2(new_n1146), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1148), .B1(new_n1158), .B2(new_n1145), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n744), .B2(new_n742), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1157), .B1(new_n1160), .B2(KEYINPUT127), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(KEYINPUT127), .B2(new_n1160), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(KEYINPUT48), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(KEYINPUT48), .B2(new_n1164), .ZN(new_n1166));
  OR3_X1    g741(.A1(new_n1157), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT46), .B1(new_n1157), .B2(G1996), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1146), .A2(new_n708), .A3(new_n712), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1167), .A2(new_n1168), .B1(new_n1145), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT47), .Z(new_n1171));
  NAND3_X1  g746(.A1(new_n1162), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1156), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g749(.A1(G227), .A2(new_n459), .ZN(new_n1176));
  NOR3_X1   g750(.A1(G229), .A2(G401), .A3(new_n1176), .ZN(new_n1177));
  AND4_X1   g751(.A1(KEYINPUT112), .A2(new_n905), .A3(new_n908), .A4(new_n909), .ZN(new_n1178));
  AOI21_X1  g752(.A(KEYINPUT112), .B1(new_n913), .B2(new_n908), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n965), .B2(new_n966), .ZN(G308));
  OAI221_X1 g755(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .C1(new_n960), .C2(new_n961), .ZN(G225));
endmodule


