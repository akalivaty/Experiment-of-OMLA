//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G50), .B(G68), .Z(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n250), .A2(G223), .B1(new_n253), .B2(G77), .ZN(new_n254));
  INV_X1    g0054(.A(G222), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n249), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n245), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n214), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n206), .B(G274), .C1(new_n259), .C2(new_n214), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n264), .A2(new_n268), .ZN(new_n270));
  INV_X1    g0070(.A(new_n214), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n206), .A2(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n263), .A2(new_n269), .B1(new_n273), .B2(G226), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n261), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G200), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(new_n261), .B2(new_n274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT66), .A2(G58), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT8), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT67), .B1(new_n284), .B2(KEYINPUT8), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n285), .A2(new_n291), .A3(KEYINPUT8), .A4(new_n286), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT64), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n296), .A3(G33), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n282), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(new_n214), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n202), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n206), .A2(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(new_n202), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT9), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n302), .A2(KEYINPUT9), .A3(new_n308), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n280), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n280), .B(new_n315), .C1(new_n311), .C2(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n309), .B1(new_n318), .B2(new_n275), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G179), .B2(new_n275), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  INV_X1    g0121(.A(G77), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n321), .B1(new_n307), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n300), .A2(KEYINPUT68), .A3(G77), .A4(new_n306), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  INV_X1    g0126(.A(new_n281), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n322), .A2(new_n213), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n297), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n301), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n304), .A2(new_n322), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT69), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n256), .A2(G232), .A3(new_n245), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n253), .A2(G107), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n260), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n263), .A2(new_n269), .B1(new_n273), .B2(G244), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G200), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT69), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n325), .A2(new_n331), .A3(new_n343), .A4(new_n332), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n334), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT70), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n334), .A2(new_n342), .A3(new_n347), .A4(new_n344), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n339), .A2(G190), .A3(new_n340), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n334), .A2(new_n344), .ZN(new_n351));
  AOI21_X1  g0151(.A(G169), .B1(new_n339), .B2(new_n340), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n339), .A2(new_n340), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n317), .A2(new_n320), .A3(new_n350), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G159), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n327), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(KEYINPUT66), .A2(G58), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT66), .A2(G58), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n216), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n359), .B1(new_n363), .B2(G20), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n253), .A2(new_n213), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n248), .A2(new_n207), .A3(new_n249), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT7), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n368), .A3(G68), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n364), .A2(new_n369), .A3(KEYINPUT16), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n301), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n253), .A2(new_n365), .A3(new_n207), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n294), .A2(new_n296), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n256), .ZN(new_n374));
  OAI211_X1 g0174(.A(G68), .B(new_n372), .C1(new_n374), .C2(new_n365), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT16), .B1(new_n375), .B2(new_n364), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n290), .A2(new_n307), .A3(new_n292), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n304), .B1(new_n290), .B2(new_n292), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT73), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n360), .A2(new_n361), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n288), .B1(new_n381), .B2(KEYINPUT8), .ZN(new_n382));
  INV_X1    g0182(.A(new_n292), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n303), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n290), .A2(new_n307), .A3(new_n292), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n371), .A2(new_n376), .B1(new_n379), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n271), .A2(new_n272), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G232), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n269), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n262), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT74), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n393), .B(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(G223), .B(new_n245), .C1(new_n251), .C2(new_n252), .ZN(new_n396));
  OAI211_X1 g0196(.A(G226), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n392), .B1(new_n260), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n260), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n263), .A2(new_n269), .B1(new_n273), .B2(G232), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n387), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT18), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n387), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n365), .B1(new_n253), .B2(new_n213), .ZN(new_n411));
  NOR4_X1   g0211(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT7), .A4(G20), .ZN(new_n412));
  INV_X1    g0212(.A(G68), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT66), .B(G58), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n201), .B1(new_n415), .B2(G68), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n416), .A2(new_n207), .B1(new_n358), .B2(new_n327), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n410), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n301), .A3(new_n370), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n401), .A2(new_n402), .A3(new_n276), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n399), .B2(G200), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT73), .B1(new_n377), .B2(new_n378), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n384), .A2(new_n380), .A3(new_n385), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n419), .A2(new_n421), .A3(new_n424), .A4(KEYINPUT17), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n407), .A2(new_n409), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n357), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n413), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n297), .B2(new_n322), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n301), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT71), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(KEYINPUT71), .A3(new_n301), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n439), .A2(KEYINPUT11), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT12), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n304), .B2(new_n413), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n303), .A2(KEYINPUT12), .A3(G68), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n442), .A2(new_n443), .B1(new_n307), .B2(new_n413), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n439), .B2(KEYINPUT11), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n273), .A2(G238), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n269), .A2(new_n388), .A3(new_n206), .A4(G274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n230), .A2(G1698), .ZN(new_n451));
  OAI221_X1 g0251(.A(new_n451), .B1(G226), .B2(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G97), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n388), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT13), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n450), .A2(new_n454), .A3(KEYINPUT13), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n447), .B(G169), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n450), .ZN(new_n459));
  INV_X1    g0259(.A(new_n454), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT13), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(G179), .A3(new_n455), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n455), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n447), .B1(new_n465), .B2(G169), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n446), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(G200), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(G190), .A3(new_n455), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n440), .A3(new_n445), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g0271(.A(new_n471), .B(KEYINPUT72), .Z(new_n472));
  NAND2_X1  g0272(.A1(new_n432), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n303), .A2(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n206), .A2(G33), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n300), .A2(new_n303), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(G97), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(KEYINPUT6), .A3(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n373), .B1(G77), .B2(new_n281), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n372), .B1(new_n374), .B2(new_n365), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n479), .B1(new_n490), .B2(new_n301), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT5), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n206), .B(G45), .C1(new_n492), .C2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n265), .A2(new_n267), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(G274), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n260), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT5), .B1(new_n265), .B2(new_n267), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(new_n388), .C1(new_n499), .C2(new_n493), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n256), .A2(G244), .A3(new_n245), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n245), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n250), .A2(G250), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n501), .B1(new_n508), .B2(new_n260), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G190), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n498), .A2(new_n500), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT76), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n498), .B2(new_n500), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n513), .A2(new_n515), .B1(new_n260), .B2(new_n508), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n491), .B(new_n510), .C1(new_n516), .C2(new_n278), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n490), .A2(new_n301), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n478), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n508), .A2(new_n260), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n318), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n501), .A2(KEYINPUT76), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n353), .B(new_n520), .C1(new_n523), .C2(new_n514), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n297), .B2(new_n481), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n256), .A2(new_n213), .A3(G68), .ZN(new_n529));
  INV_X1    g0329(.A(new_n453), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n373), .B1(KEYINPUT19), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n528), .B(new_n529), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n301), .B1(new_n304), .B2(new_n329), .ZN(new_n534));
  INV_X1    g0334(.A(new_n329), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n477), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n206), .A2(new_n496), .A3(G45), .ZN(new_n539));
  INV_X1    g0339(.A(G250), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n268), .B2(G1), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n388), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n256), .A2(G238), .A3(new_n245), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n256), .A2(G244), .A3(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n260), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n353), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G169), .B2(new_n548), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(G190), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n477), .A2(G87), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n534), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n548), .A2(new_n278), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n538), .A2(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT77), .B1(new_n526), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n551), .A2(new_n534), .A3(new_n552), .ZN(new_n557));
  INV_X1    g0357(.A(new_n554), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n548), .A2(G169), .ZN(new_n559));
  AOI211_X1 g0359(.A(G179), .B(new_n543), .C1(new_n547), .C2(new_n260), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n557), .A2(new_n558), .B1(new_n561), .B2(new_n537), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n517), .A3(new_n563), .A4(new_n525), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n256), .A2(new_n213), .A3(G87), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT79), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(KEYINPUT24), .B1(KEYINPUT23), .B2(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(G20), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(KEYINPUT23), .A2(G107), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n373), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n567), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n569), .B1(new_n567), .B2(new_n574), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n301), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n477), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n303), .A2(G107), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT80), .B(KEYINPUT25), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G294), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n257), .C2(new_n540), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n260), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(new_n388), .C1(new_n499), .C2(new_n493), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n498), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n589), .A2(new_n276), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(G200), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n578), .A2(new_n583), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(G169), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT81), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n587), .A2(new_n588), .A3(G179), .A4(new_n498), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(new_n596), .A3(G169), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n583), .ZN(new_n599));
  INV_X1    g0399(.A(new_n577), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n575), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n599), .B1(new_n601), .B2(new_n301), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n592), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G116), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n299), .A2(new_n214), .B1(G20), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n506), .B1(new_n481), .B2(G33), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n373), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n605), .B(KEYINPUT20), .C1(new_n373), .C2(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n303), .A2(G116), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n477), .B2(G116), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT78), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT78), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(G270), .B(new_n388), .C1(new_n499), .C2(new_n493), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n498), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n250), .A2(G264), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n256), .A2(G257), .A3(new_n245), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n253), .A2(G303), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n260), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G190), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n626), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n619), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n318), .B1(new_n621), .B2(new_n626), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT78), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT78), .B1(new_n611), .B2(new_n613), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n627), .B(G179), .C1(new_n633), .C2(new_n634), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n632), .B(KEYINPUT21), .C1(new_n633), .C2(new_n634), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n631), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n603), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n474), .A2(new_n565), .A3(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n427), .A2(new_n428), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n356), .A2(KEYINPUT83), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT83), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n351), .A2(new_n355), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n470), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n643), .B1(new_n647), .B2(new_n467), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n407), .A2(new_n409), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n317), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n538), .A2(new_n550), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n562), .A2(new_n652), .A3(KEYINPUT26), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n555), .B2(new_n525), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n597), .A2(new_n595), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n594), .B1(new_n578), .B2(new_n583), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT82), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n638), .A2(new_n639), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT21), .B1(new_n618), .B2(new_n632), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n637), .A2(KEYINPUT82), .A3(new_n638), .A4(new_n639), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n592), .A2(new_n562), .A3(new_n525), .A4(new_n517), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n656), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n320), .B(new_n650), .C1(new_n473), .C2(new_n667), .ZN(G369));
  INV_X1    g0468(.A(new_n603), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n206), .A2(G13), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT27), .B1(new_n373), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT27), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n213), .A2(new_n672), .A3(new_n206), .A4(G13), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n673), .A3(G213), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT84), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G343), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n669), .B1(new_n602), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n658), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT87), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n619), .A2(new_n678), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n640), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n662), .A2(new_n663), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n689), .B2(new_n686), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT85), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT85), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n692), .B(new_n687), .C1(new_n689), .C2(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(KEYINPUT86), .B(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n684), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  AOI211_X1 g0497(.A(KEYINPUT87), .B(new_n695), .C1(new_n691), .C2(new_n693), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n683), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n660), .A2(new_n661), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n680), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n669), .A2(new_n701), .B1(new_n658), .B2(new_n678), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n210), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n494), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n206), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n532), .A2(new_n604), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n706), .A2(new_n708), .B1(new_n218), .B2(new_n705), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n666), .A2(new_n711), .A3(new_n678), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT88), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n526), .B(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n658), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n700), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n562), .A3(new_n592), .A4(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n680), .B1(new_n717), .B2(new_n656), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n712), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n565), .A2(new_n641), .A3(new_n678), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n627), .A2(G179), .A3(new_n548), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n520), .B1(new_n523), .B2(new_n514), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n589), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n629), .A2(new_n353), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n548), .A2(new_n588), .A3(new_n587), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(new_n509), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n725), .A4(new_n509), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n680), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n720), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n719), .B1(new_n696), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n710), .B1(new_n735), .B2(G1), .ZN(G364));
  AOI21_X1  g0536(.A(new_n214), .B1(G20), .B2(new_n318), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n213), .A2(new_n353), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G190), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n278), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n373), .A2(new_n276), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n741), .A2(G311), .B1(G283), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G294), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n276), .A2(G200), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n213), .B1(new_n353), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n738), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(G190), .A3(new_n278), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n750), .A2(new_n276), .A3(new_n278), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G326), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n738), .A2(new_n747), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G322), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n742), .A2(G20), .A3(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n256), .B1(new_n760), .B2(G303), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n753), .A2(new_n755), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n213), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n749), .B(new_n762), .C1(G329), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n743), .A2(new_n482), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n253), .B(new_n769), .C1(G87), .C2(new_n760), .ZN(new_n770));
  INV_X1    g0570(.A(new_n754), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n202), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n763), .A2(G159), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n751), .A2(G68), .B1(new_n773), .B2(KEYINPUT32), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(KEYINPUT32), .B2(new_n773), .ZN(new_n775));
  INV_X1    g0575(.A(new_n748), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G97), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n777), .B1(new_n756), .B2(new_n381), .C1(new_n322), .C2(new_n740), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n772), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n737), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n213), .A2(G13), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT89), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G45), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n706), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n704), .A2(new_n253), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G355), .B1(new_n604), .B2(new_n704), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n704), .A2(new_n256), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G45), .B2(new_n217), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n240), .A2(new_n268), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT90), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n737), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n791), .B2(new_n792), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n780), .B(new_n785), .C1(new_n793), .C2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT92), .Z(new_n800));
  INV_X1    g0600(.A(new_n796), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n694), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n694), .A2(new_n696), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n698), .A2(new_n697), .A3(new_n804), .A4(new_n785), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n803), .A2(new_n805), .ZN(G396));
  INV_X1    g0606(.A(new_n737), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n795), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G143), .A2(new_n757), .B1(new_n741), .B2(G159), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n751), .A2(G150), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n771), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n744), .A2(G68), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n253), .B1(new_n760), .B2(G50), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n381), .C2(new_n748), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n767), .B2(G132), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n256), .B1(new_n760), .B2(G107), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n777), .B(new_n818), .C1(new_n771), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G283), .B2(new_n751), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n744), .A2(G87), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n757), .B2(G294), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n604), .B2(new_n740), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G311), .B2(new_n767), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n813), .A2(new_n817), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n785), .B1(G77), .B2(new_n808), .C1(new_n826), .C2(new_n807), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n350), .A2(KEYINPUT94), .A3(new_n356), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n351), .A2(new_n680), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT94), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n350), .A2(new_n831), .A3(new_n356), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n829), .B1(new_n644), .B2(new_n646), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n827), .B1(new_n794), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n667), .B2(new_n680), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n832), .A2(new_n833), .B1(new_n828), .B2(new_n829), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n666), .A2(new_n678), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n734), .A2(new_n696), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n785), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n836), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  OR2_X1    g0645(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(G116), .A3(new_n215), .A4(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(KEYINPUT95), .B(KEYINPUT36), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n218), .A2(G77), .A3(new_n362), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n851), .A2(KEYINPUT96), .B1(G50), .B2(new_n413), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(KEYINPUT96), .B2(new_n851), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n206), .A2(G13), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n364), .B2(new_n369), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n371), .A2(new_n855), .B1(new_n379), .B2(new_n386), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n676), .A2(new_n677), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n429), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n405), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n859), .A3(new_n425), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n387), .A2(new_n858), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n406), .A2(new_n865), .A3(new_n866), .A4(new_n425), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n868), .A3(KEYINPUT38), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n861), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n356), .A2(new_n680), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n839), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n678), .B1(new_n440), .B2(new_n445), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n467), .A2(new_n470), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT97), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n876), .B(new_n879), .C1(new_n464), .C2(new_n466), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n876), .B1(new_n464), .B2(new_n466), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT97), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n872), .B1(new_n884), .B2(KEYINPUT98), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT98), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n875), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n649), .A2(new_n857), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n467), .A2(new_n680), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n419), .A2(new_n421), .A3(new_n424), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n419), .A2(new_n424), .B1(new_n404), .B2(new_n400), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n866), .B1(new_n894), .B2(new_n865), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n896));
  INV_X1    g0696(.A(new_n865), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n895), .A2(new_n896), .B1(new_n429), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n406), .A2(new_n865), .A3(new_n425), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(KEYINPUT99), .A3(new_n867), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n869), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT100), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n429), .A2(new_n860), .B1(new_n864), .B2(new_n867), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT39), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n429), .A2(new_n897), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT99), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n899), .A2(new_n909), .A3(KEYINPUT37), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n901), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT100), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n870), .B2(new_n871), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n905), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT101), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT101), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n905), .A2(new_n915), .A3(new_n916), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n891), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n890), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n650), .A2(new_n320), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n719), .B2(new_n474), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT102), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n883), .A2(new_n830), .A3(new_n834), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n734), .A2(KEYINPUT40), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n902), .A2(new_n870), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n883), .A2(new_n830), .A3(new_n834), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n720), .B2(new_n733), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n913), .A2(new_n869), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n932), .A2(KEYINPUT102), .A3(KEYINPUT40), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n870), .B2(new_n871), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n474), .A2(new_n734), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n695), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n925), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n206), .B2(new_n782), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n925), .A2(new_n942), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n850), .B1(new_n853), .B2(new_n854), .C1(new_n944), .C2(new_n945), .ZN(G367));
  INV_X1    g0746(.A(new_n788), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n797), .B1(new_n210), .B2(new_n329), .C1(new_n947), .C2(new_n236), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n785), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n534), .A2(new_n552), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n680), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n562), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n651), .A2(new_n950), .A3(new_n680), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n754), .A2(G143), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n253), .B1(new_n760), .B2(new_n415), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(new_n322), .C2(new_n743), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G50), .A2(new_n741), .B1(new_n757), .B2(G150), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n776), .A2(G68), .ZN(new_n959));
  INV_X1    g0759(.A(new_n763), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n959), .C1(new_n811), .C2(new_n960), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n957), .B(new_n961), .C1(G159), .C2(new_n751), .ZN(new_n962));
  INV_X1    g0762(.A(new_n751), .ZN(new_n963));
  INV_X1    g0763(.A(G311), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n746), .A2(new_n963), .B1(new_n771), .B2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n741), .A2(G283), .B1(G97), .B2(new_n744), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n482), .B2(new_n748), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n760), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT46), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n759), .B2(new_n604), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n253), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n763), .A2(G317), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n819), .B2(new_n756), .ZN(new_n973));
  NOR4_X1   g0773(.A1(new_n965), .A2(new_n967), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n962), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n949), .B1(new_n801), .B2(new_n954), .C1(new_n976), .C2(new_n807), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n783), .A2(G1), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT105), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n735), .ZN(new_n982));
  INV_X1    g0782(.A(new_n697), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n694), .A2(new_n684), .A3(new_n696), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n669), .A2(new_n701), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n682), .B1(new_n700), .B2(new_n680), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n697), .B2(new_n698), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n519), .A2(new_n680), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n714), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n652), .A2(new_n680), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n702), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(KEYINPUT44), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n994), .A2(new_n702), .A3(new_n997), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n994), .A2(KEYINPUT45), .A3(new_n702), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT45), .B1(new_n994), .B2(new_n702), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n996), .A2(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(new_n683), .C1(new_n698), .C2(new_n697), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n990), .A2(new_n1002), .A3(new_n735), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT104), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n699), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1001), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(KEYINPUT104), .A3(new_n699), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n982), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n705), .B(KEYINPUT41), .Z(new_n1011));
  OAI21_X1  g0811(.A(new_n981), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n985), .B1(new_n992), .B2(new_n993), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT42), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT43), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n954), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n525), .B1(new_n992), .B2(new_n715), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n678), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n954), .B(new_n1015), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(KEYINPUT103), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT103), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1005), .A2(new_n994), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1023), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n978), .B1(new_n1012), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(G387));
  NAND2_X1  g0828(.A1(new_n990), .A2(new_n735), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n982), .A2(new_n987), .A3(new_n989), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n705), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n682), .A2(new_n796), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n786), .A2(new_n707), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(G107), .B2(new_n210), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n233), .A2(new_n268), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT106), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n326), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n947), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n797), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n785), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT107), .B(G150), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n960), .A2(new_n1044), .B1(new_n202), .B2(new_n756), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n740), .A2(new_n413), .B1(new_n748), .B2(new_n329), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n754), .A2(G159), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n293), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n751), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n256), .B1(new_n759), .B2(new_n322), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n744), .B2(G97), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n256), .B1(new_n763), .B2(G326), .ZN(new_n1054));
  INV_X1    g0854(.A(G283), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n748), .A2(new_n1055), .B1(new_n746), .B2(new_n759), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G303), .A2(new_n741), .B1(new_n757), .B2(G317), .ZN(new_n1057));
  INV_X1    g0857(.A(G322), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1057), .B1(new_n963), .B2(new_n964), .C1(new_n1058), .C2(new_n771), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1054), .B1(new_n604), .B2(new_n743), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1053), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1043), .B1(new_n1066), .B2(new_n737), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n990), .A2(new_n980), .B1(new_n1032), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1031), .A2(new_n1068), .ZN(G393));
  XNOR2_X1  g0869(.A(new_n1002), .B(KEYINPUT108), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n992), .A2(new_n796), .A3(new_n993), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n797), .B1(new_n481), .B2(new_n210), .C1(new_n947), .C2(new_n243), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n785), .A2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n754), .A2(G317), .B1(G311), .B2(new_n757), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n960), .A2(new_n1058), .B1(new_n604), .B2(new_n748), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G294), .B2(new_n741), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n253), .B1(new_n759), .B2(new_n1055), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n769), .B(new_n1080), .C1(new_n751), .C2(G303), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n754), .A2(G150), .B1(G159), .B2(new_n757), .ZN(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n763), .A2(G143), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n413), .B2(new_n759), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n253), .B(new_n822), .C1(new_n1087), .C2(KEYINPUT110), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(KEYINPUT110), .C2(new_n1087), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n776), .A2(G77), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n326), .B2(new_n740), .C1(new_n963), .C2(new_n202), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT111), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1082), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1074), .B1(new_n1093), .B2(new_n737), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1071), .A2(new_n980), .B1(new_n1072), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n990), .A2(new_n1002), .A3(new_n735), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n705), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1029), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1071), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1095), .B1(new_n1099), .B2(new_n1101), .ZN(G390));
  NAND4_X1  g0902(.A1(new_n734), .A2(new_n432), .A3(G330), .A4(new_n472), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT115), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n924), .ZN(new_n1105));
  INV_X1    g0905(.A(G330), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1106), .B(new_n835), .C1(new_n720), .C2(new_n733), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n883), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n841), .A2(new_n835), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n883), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n875), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n734), .A2(new_n696), .A3(new_n838), .A4(new_n883), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT114), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n873), .B1(new_n718), .B2(new_n838), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1107), .A2(new_n883), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1105), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n884), .A2(new_n891), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n918), .A2(new_n920), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n883), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n891), .B(new_n933), .C1(new_n1114), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT113), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1108), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n1122), .A3(new_n1113), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT113), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(new_n1127), .A3(new_n1126), .A4(new_n1117), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n705), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1132), .A2(new_n980), .A3(new_n1127), .A4(new_n1126), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n918), .A2(new_n794), .A3(new_n920), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1090), .B1(new_n756), .B2(new_n604), .C1(new_n481), .C2(new_n740), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n256), .B1(new_n760), .B2(G87), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n814), .A2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n963), .B2(new_n482), .C1(new_n1055), .C2(new_n771), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(G294), .C2(new_n767), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n256), .B1(new_n202), .B2(new_n743), .C1(new_n766), .C2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT117), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n757), .A2(G132), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G128), .A2(new_n754), .B1(new_n751), .B2(G137), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n759), .A2(new_n1044), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT116), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1150), .A2(new_n741), .B1(G159), .B2(new_n776), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1141), .B1(new_n1144), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n785), .B1(new_n1049), .B2(new_n808), .C1(new_n1153), .C2(new_n807), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT118), .Z(new_n1155));
  NAND2_X1  g0955(.A1(new_n1136), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1135), .A2(new_n1156), .A3(KEYINPUT119), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT119), .B1(new_n1135), .B2(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1134), .B1(new_n1157), .B2(new_n1158), .ZN(G378));
  AOI22_X1  g0959(.A1(new_n930), .A2(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n317), .A2(new_n320), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n309), .A2(new_n857), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1160), .A2(G330), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1160), .B2(G330), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n921), .B2(new_n890), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1165), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n939), .B2(new_n1106), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n921), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n885), .A2(new_n887), .B1(new_n649), .B2(new_n857), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1160), .A2(G330), .A3(new_n1165), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n794), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n785), .B1(G50), .B2(new_n808), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n256), .A2(new_n494), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G50), .B(new_n1178), .C1(new_n247), .C2(new_n264), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n256), .B(new_n494), .C1(new_n760), .C2(G77), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n959), .B(new_n1180), .C1(new_n771), .C2(new_n604), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G97), .B2(new_n751), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n743), .A2(new_n381), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n756), .A2(new_n482), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n535), .C2(new_n741), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1182), .B(new_n1185), .C1(new_n1055), .C2(new_n766), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1179), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n763), .A2(G124), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(G41), .C1(new_n744), .C2(G159), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1150), .A2(new_n760), .B1(new_n776), .B2(G150), .ZN(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n756), .C1(new_n771), .C2(new_n1142), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n751), .A2(G132), .B1(G137), .B2(new_n741), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT59), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1189), .B(new_n1190), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1177), .B1(new_n1201), .B2(new_n737), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1175), .A2(new_n980), .B1(new_n1176), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  AOI211_X1 g1004(.A(KEYINPUT113), .B(new_n1108), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1127), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1129), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1105), .B1(new_n1207), .B2(new_n1117), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1105), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1133), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(KEYINPUT121), .A3(new_n1210), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1133), .A2(new_n1213), .B1(new_n1174), .B2(new_n1168), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n705), .B1(new_n1217), .B2(KEYINPUT57), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1203), .B1(new_n1216), .B2(new_n1218), .ZN(G375));
  NAND2_X1  g1019(.A1(new_n1116), .A2(new_n1111), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1121), .A2(new_n794), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n785), .B1(G68), .B2(new_n808), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  INV_X1    g1023(.A(G132), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n771), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n754), .A2(KEYINPUT122), .A3(G132), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n1192), .C2(new_n766), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n253), .B(new_n1183), .C1(G159), .C2(new_n760), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n741), .A2(G150), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n757), .A2(G137), .B1(new_n776), .B2(G50), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n751), .A2(new_n1150), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n253), .B1(new_n759), .B2(new_n481), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n744), .B2(G77), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n963), .B2(new_n604), .C1(new_n746), .C2(new_n771), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n757), .A2(G283), .B1(new_n776), .B2(new_n535), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n482), .B2(new_n740), .C1(new_n766), .C2(new_n819), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1227), .A2(new_n1232), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1222), .B1(new_n1238), .B2(new_n737), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1220), .A2(new_n980), .B1(new_n1221), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1011), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1118), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1220), .A2(new_n1213), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(G381));
  NOR2_X1   g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1203), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1214), .A2(KEYINPUT121), .A3(new_n1210), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT121), .B1(new_n1214), .B2(new_n1210), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1217), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1098), .B1(new_n1253), .B2(new_n1209), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1249), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1247), .A2(new_n1027), .A3(new_n1248), .A4(new_n1255), .ZN(G407));
  INV_X1    g1056(.A(G343), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1248), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G407), .A2(G213), .A3(new_n1260), .ZN(G409));
  OAI211_X1 g1061(.A(G378), .B(new_n1203), .C1(new_n1216), .C2(new_n1218), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1217), .A2(new_n1241), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1203), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1248), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1220), .A2(new_n1213), .A3(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(new_n1098), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1117), .A2(new_n1267), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1243), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1240), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n844), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(G384), .A3(new_n1240), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1266), .A2(new_n1258), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1259), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1275), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1259), .A2(G2897), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1273), .A2(new_n1274), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G378), .B1(new_n1203), .B2(new_n1263), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1255), .B2(G378), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1288), .B2(new_n1259), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1277), .A2(new_n1278), .A3(new_n1281), .A4(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1291), .A2(new_n1245), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1292), .B1(new_n1027), .B2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1291), .A2(new_n1245), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1023), .B(new_n1024), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1241), .B1(new_n1097), .B2(new_n982), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n981), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1295), .B1(new_n1298), .B2(new_n978), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1294), .A2(G390), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G390), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1290), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(KEYINPUT123), .B(new_n1286), .C1(new_n1288), .C2(new_n1259), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT123), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1285), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1283), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1279), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1278), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1276), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT125), .B1(new_n1276), .B2(new_n1311), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1279), .A2(new_n1314), .A3(KEYINPUT63), .A4(new_n1275), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1309), .A2(new_n1312), .A3(new_n1313), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1303), .A2(new_n1316), .ZN(G405));
  NAND2_X1  g1117(.A1(G375), .A2(new_n1248), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1262), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1275), .A2(KEYINPUT126), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1318), .A2(new_n1262), .A3(new_n1320), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1325), .A2(new_n1326), .B1(new_n1327), .B2(new_n1302), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1327), .B2(new_n1302), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1302), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1325), .A2(new_n1330), .A3(KEYINPUT127), .A4(new_n1326), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(G402));
endmodule


