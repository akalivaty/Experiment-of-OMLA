//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n459), .A2(new_n460), .A3(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n460), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n463), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(G2104), .B2(new_n465), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n462), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(G2105), .A2(new_n474), .B1(new_n478), .B2(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n469), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n466), .A2(new_n461), .A3(G2105), .A4(new_n463), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT69), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n484), .B(new_n488), .C1(G136), .C2(new_n468), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n466), .A2(new_n461), .A3(new_n463), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n472), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n509), .A2(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n505), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n509), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n520), .B(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n504), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n509), .A2(new_n532), .B1(new_n515), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  NOR2_X1   g110(.A1(new_n512), .A2(new_n511), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  INV_X1    g112(.A(G68), .ZN(new_n538));
  INV_X1    g113(.A(G543), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n542), .B1(new_n538), .B2(new_n539), .C1(new_n536), .C2(new_n537), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(G651), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n539), .B1(new_n506), .B2(new_n507), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n519), .A2(G81), .B1(G43), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(G860), .A3(new_n546), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n508), .A2(new_n502), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(G91), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n545), .A2(new_n556), .A3(G53), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n536), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n555), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  OR2_X1    g143(.A1(new_n505), .A2(new_n517), .ZN(G303));
  NAND3_X1  g144(.A1(new_n552), .A2(G87), .A3(new_n554), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n536), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n545), .B2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n536), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G48), .B2(new_n545), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n552), .A2(G86), .A3(new_n554), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n504), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n509), .A2(new_n583), .B1(new_n515), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n552), .A2(G92), .A3(new_n554), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n590), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n552), .A2(G92), .A3(new_n554), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n536), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n545), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n544), .A2(new_n546), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n599), .A2(new_n606), .ZN(new_n609));
  MUX2_X1   g184(.A(new_n608), .B(new_n609), .S(G868), .Z(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n478), .A2(new_n493), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  XOR2_X1   g188(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n613), .B(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n618));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n485), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n468), .B2(G135), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2096), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n623), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT77), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n629), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT78), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT80), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G1986), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT79), .ZN(new_n672));
  INV_X1    g247(.A(G1981), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT79), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n673), .B1(new_n672), .B2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n659), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(G1986), .A3(new_n676), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n658), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n681), .A3(new_n658), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n684), .ZN(new_n687));
  INV_X1    g262(.A(new_n685), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n682), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(G229));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G6), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(G23), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G288), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n694), .A2(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n692), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G1971), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(G1971), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n703), .B(new_n704), .C1(new_n694), .C2(new_n695), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT34), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n692), .A2(G24), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n586), .B2(new_n692), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT83), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(new_n659), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT81), .B(G29), .Z(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n716));
  INV_X1    g291(.A(G119), .ZN(new_n717));
  INV_X1    g292(.A(G131), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n716), .B1(new_n717), .B2(new_n485), .C1(new_n467), .C2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT82), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT82), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n713), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n714), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n712), .A2(KEYINPUT84), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n708), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT85), .B(KEYINPUT36), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n723), .A2(G35), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G162), .B2(new_n723), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT29), .Z(new_n734));
  INV_X1    g309(.A(G2090), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n692), .A2(G21), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G168), .B2(new_n692), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT92), .Z(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT25), .Z(new_n745));
  INV_X1    g320(.A(G139), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n467), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  INV_X1    g323(.A(G127), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n472), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n465), .B1(new_n750), .B2(KEYINPUT88), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(KEYINPUT88), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n743), .B1(new_n753), .B2(new_n742), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G2072), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT90), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  INV_X1    g333(.A(G129), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n485), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n478), .A2(G105), .ZN(new_n761));
  INV_X1    g336(.A(G141), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n467), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n742), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n742), .B2(G32), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT27), .B(G1996), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT91), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n766), .A2(new_n768), .B1(G2072), .B2(new_n754), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n755), .B(new_n769), .C1(new_n768), .C2(new_n766), .ZN(new_n770));
  MUX2_X1   g345(.A(G19), .B(new_n608), .S(G16), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1341), .ZN(new_n772));
  INV_X1    g347(.A(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT30), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n692), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n692), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n778), .B1(new_n780), .B2(G1961), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G34), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n713), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT89), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n480), .B2(new_n742), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n780), .A2(G1961), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n622), .B2(new_n713), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n772), .A2(new_n781), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n737), .A2(new_n741), .A3(new_n770), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n740), .A2(G1966), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT93), .Z(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(KEYINPUT94), .B2(new_n736), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n713), .A2(G26), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n468), .A2(G140), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT86), .ZN(new_n798));
  INV_X1    g373(.A(G128), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n485), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT87), .ZN(new_n801));
  OR2_X1    g376(.A1(G104), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n796), .B1(new_n805), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2067), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n692), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n599), .B2(new_n692), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1348), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n723), .A2(G27), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n723), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2078), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n692), .A2(G20), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT23), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n565), .B2(new_n692), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1956), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n810), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n807), .B(new_n818), .C1(new_n734), .C2(new_n735), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n791), .A2(new_n794), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n731), .A2(new_n820), .ZN(G311));
  NAND2_X1  g396(.A1(new_n731), .A2(new_n820), .ZN(G150));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT96), .B(G55), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n545), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n508), .A2(new_n502), .A3(G93), .ZN(new_n826));
  OAI21_X1  g401(.A(G67), .B1(new_n512), .B2(new_n511), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n504), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n825), .B(new_n826), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n832), .A2(KEYINPUT95), .A3(new_n504), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n823), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n825), .A2(new_n826), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT95), .B1(new_n832), .B2(new_n504), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n829), .A2(new_n830), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT97), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n599), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n834), .A2(new_n608), .A3(new_n838), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n544), .B(new_n546), .C1(new_n831), .C2(new_n833), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n843), .B(new_n846), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n841), .B1(new_n849), .B2(new_n851), .ZN(G145));
  XOR2_X1   g427(.A(KEYINPUT99), .B(G37), .Z(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n720), .A2(KEYINPUT98), .A3(new_n721), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT98), .B1(new_n720), .B2(new_n721), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n613), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(new_n613), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n855), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n764), .B(new_n753), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n858), .B2(new_n861), .ZN(new_n865));
  OR2_X1    g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n867));
  INV_X1    g442(.A(G130), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n485), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n468), .B2(G142), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(G164), .B1(new_n798), .B2(new_n804), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n798), .A2(new_n804), .A3(G164), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n873), .A2(new_n871), .A3(new_n874), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n864), .A2(new_n865), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n865), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n863), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n480), .B(new_n621), .ZN(new_n882));
  XNOR2_X1  g457(.A(G162), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n877), .A2(new_n880), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n854), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(G395));
  NAND2_X1  g464(.A1(new_n691), .A2(G166), .ZN(new_n890));
  NAND2_X1  g465(.A1(G303), .A2(G305), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n896));
  NAND2_X1  g471(.A1(G288), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n570), .A2(KEYINPUT101), .A3(new_n573), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(G290), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G290), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n893), .B(new_n895), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n903), .A2(KEYINPUT102), .A3(new_n892), .A4(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT42), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n598), .A2(new_n565), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n598), .A2(new_n565), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n598), .A2(new_n912), .A3(new_n565), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n598), .B2(new_n565), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(new_n914), .A3(new_n907), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n911), .B1(new_n915), .B2(KEYINPUT41), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n846), .B(new_n609), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n907), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n910), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n906), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n906), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n839), .A2(new_n602), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n928));
  XNOR2_X1  g503(.A(G331), .B(new_n928), .ZN(G295));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(KEYINPUT104), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n531), .B2(new_n534), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n844), .A2(new_n934), .A3(new_n845), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n844), .B2(new_n845), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n936), .A2(new_n937), .A3(G286), .ZN(new_n938));
  INV_X1    g513(.A(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n846), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G168), .B1(new_n940), .B2(new_n935), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n916), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n902), .A2(new_n904), .ZN(new_n943));
  OAI21_X1  g518(.A(G286), .B1(new_n936), .B2(new_n937), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(G168), .A3(new_n935), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n945), .A3(new_n920), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT105), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n942), .A2(new_n949), .A3(new_n943), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n943), .B1(new_n942), .B2(new_n946), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(new_n953), .A3(G37), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n920), .A2(new_n956), .A3(new_n908), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n913), .A2(new_n914), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n909), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n920), .B2(new_n908), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(new_n938), .B2(new_n941), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n946), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n854), .B1(new_n963), .B2(new_n905), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n951), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n930), .B(new_n955), .C1(new_n966), .C2(KEYINPUT43), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n952), .A2(KEYINPUT43), .A3(G37), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n951), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT44), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n953), .B1(new_n951), .B2(new_n964), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n930), .B1(new_n951), .B2(new_n968), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT107), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n967), .B1(new_n973), .B2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n495), .B2(new_n499), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n469), .A2(new_n479), .A3(G40), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1996), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT108), .Z(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  INV_X1    g562(.A(new_n764), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n985), .B(KEYINPUT108), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT109), .B1(new_n990), .B2(new_n764), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n720), .A2(new_n725), .A3(new_n721), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n725), .B1(new_n720), .B2(new_n721), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n983), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n805), .B(G2067), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n764), .A2(new_n984), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n983), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n992), .A2(KEYINPUT127), .A3(new_n995), .A4(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n995), .B(new_n998), .C1(new_n989), .C2(new_n991), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT127), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G290), .A2(G1986), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n983), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n999), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n993), .B(new_n998), .C1(new_n989), .C2(new_n991), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(G2067), .B2(new_n805), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n983), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n996), .A2(new_n988), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n983), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT126), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n990), .B2(KEYINPUT46), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n986), .A2(KEYINPUT126), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1012), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT47), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1012), .B(new_n1019), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1006), .A2(new_n1009), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n982), .B2(new_n979), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G86), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n578), .B1(new_n1025), .B2(new_n515), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G1981), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT112), .B(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n578), .A2(new_n579), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI211_X1 g609(.A(KEYINPUT114), .B(new_n1031), .C1(new_n1027), .C2(new_n1029), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1024), .B(new_n1030), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G288), .A2(G1976), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1036), .A2(new_n1037), .B1(new_n691), .B2(new_n1028), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n500), .A2(new_n1039), .A3(new_n978), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n469), .A2(new_n479), .A3(G40), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT110), .B(G2090), .ZN(new_n1044));
  INV_X1    g619(.A(G1971), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT45), .B(new_n978), .C1(new_n495), .C2(new_n499), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1046), .A3(new_n981), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1043), .A2(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G303), .A2(G8), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT55), .ZN(new_n1051));
  OR3_X1    g626(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n570), .A2(KEYINPUT111), .A3(new_n573), .A4(G1976), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1024), .A2(new_n1053), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1053), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT52), .B1(new_n1023), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1036), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g636(.A1(new_n1038), .A2(new_n1023), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1036), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1047), .A2(new_n1045), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1044), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1051), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1046), .A2(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1046), .A2(KEYINPUT115), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1041), .A3(new_n981), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1966), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(new_n1073), .B1(new_n1043), .B2(new_n786), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1074), .A2(new_n1049), .A3(G286), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1063), .A2(new_n1069), .A3(new_n1052), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1068), .A2(KEYINPUT116), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1067), .A2(new_n1080), .A3(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1051), .A3(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1061), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1082), .A2(new_n1084), .A3(KEYINPUT63), .A4(new_n1075), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1062), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G168), .A2(new_n1049), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT123), .B1(new_n1074), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1043), .A2(new_n786), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1087), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(KEYINPUT51), .B(new_n1088), .C1(new_n1074), .C2(new_n1049), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(G8), .C1(new_n1092), .C2(G286), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT62), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1063), .A2(new_n1069), .A3(new_n1052), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1065), .A2(KEYINPUT119), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1040), .A2(new_n1041), .A3(new_n1104), .A4(new_n1042), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1047), .B2(G2078), .ZN(new_n1108));
  INV_X1    g683(.A(G2078), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT53), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1106), .B(new_n1108), .C1(new_n1110), .C2(new_n1072), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1095), .A2(new_n1114), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1100), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1086), .A2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n981), .A2(new_n1046), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1041), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1956), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1065), .A2(KEYINPUT117), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT117), .B1(new_n1065), .B2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n555), .A2(new_n564), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(KEYINPUT118), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G299), .B(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1128), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(new_n1120), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT61), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n982), .B2(new_n979), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1047), .B2(G1996), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n608), .A2(KEYINPUT122), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT59), .Z(new_n1138));
  NOR2_X1   g713(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1348), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1102), .A2(new_n1140), .A3(new_n1105), .ZN(new_n1141));
  OR3_X1    g716(.A1(new_n982), .A2(G2067), .A3(new_n979), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(KEYINPUT120), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT120), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT60), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1143), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1151), .A3(new_n599), .ZN(new_n1152));
  OAI211_X1 g727(.A(KEYINPUT60), .B(new_n598), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1129), .A2(new_n1131), .A3(KEYINPUT61), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1139), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1144), .A2(new_n1145), .A3(new_n598), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1129), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1156), .B(new_n1131), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1131), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT121), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1155), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1110), .B1(new_n1041), .B2(KEYINPUT125), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1164), .B(new_n1118), .C1(KEYINPUT125), .C2(new_n1041), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1106), .A2(new_n1108), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1166), .B2(G171), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(G171), .B2(new_n1111), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1112), .B1(G171), .B2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1163), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1101), .ZN(new_n1171));
  AND4_X1   g746(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1099), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1117), .B1(new_n1162), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n586), .A2(new_n659), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n983), .B1(new_n1003), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n992), .A2(new_n1175), .A3(new_n995), .A4(new_n998), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1022), .B1(new_n1173), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g752(.A(new_n955), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n1179));
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  NOR3_X1   g754(.A1(G401), .A2(new_n1180), .A3(G227), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n686), .A2(new_n689), .A3(new_n1181), .ZN(new_n1182));
  NOR3_X1   g756(.A1(new_n1179), .A2(new_n887), .A3(new_n1182), .ZN(G308));
  NOR2_X1   g757(.A1(new_n887), .A2(new_n1182), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n1184), .B(new_n955), .C1(KEYINPUT43), .C2(new_n966), .ZN(G225));
endmodule


