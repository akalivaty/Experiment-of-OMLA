

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XNOR2_X1 U324 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U325 ( .A(n423), .B(KEYINPUT31), .Z(n292) );
  NAND2_X1 U326 ( .A1(n513), .A2(n521), .ZN(n465) );
  INV_X1 U327 ( .A(KEYINPUT25), .ZN(n467) );
  XNOR2_X1 U328 ( .A(n468), .B(n467), .ZN(n474) );
  XNOR2_X1 U329 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n398) );
  INV_X1 U330 ( .A(KEYINPUT54), .ZN(n412) );
  XNOR2_X1 U331 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U332 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U333 ( .A(n412), .B(KEYINPUT118), .ZN(n413) );
  XNOR2_X1 U334 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n479) );
  XNOR2_X1 U335 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U336 ( .A(n480), .B(n479), .ZN(n497) );
  XNOR2_X1 U337 ( .A(n581), .B(KEYINPUT41), .ZN(n552) );
  INV_X1 U338 ( .A(n552), .ZN(n567) );
  XNOR2_X1 U339 ( .A(n410), .B(n409), .ZN(n513) );
  XNOR2_X1 U340 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U341 ( .A(G92GAT), .B(KEYINPUT106), .ZN(n482) );
  XNOR2_X1 U342 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n483), .B(n482), .ZN(G1337GAT) );
  XNOR2_X1 U344 ( .A(KEYINPUT2), .B(KEYINPUT87), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n293), .B(KEYINPUT3), .ZN(n294) );
  XOR2_X1 U346 ( .A(n294), .B(KEYINPUT88), .Z(n296) );
  XNOR2_X1 U347 ( .A(G141GAT), .B(G155GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n428) );
  XOR2_X1 U349 ( .A(G127GAT), .B(KEYINPUT0), .Z(n298) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(KEYINPUT81), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n445) );
  XOR2_X1 U352 ( .A(G162GAT), .B(n445), .Z(n300) );
  XOR2_X1 U353 ( .A(G113GAT), .B(G1GAT), .Z(n319) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(n319), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n428), .B(n301), .ZN(n314) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(G85GAT), .Z(n303) );
  XNOR2_X1 U358 ( .A(G120GAT), .B(G148GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n305) );
  XNOR2_X1 U361 ( .A(KEYINPUT91), .B(G57GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n312) );
  XOR2_X1 U364 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n309) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U367 ( .A(KEYINPUT6), .B(n310), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n529) );
  XOR2_X1 U370 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n316) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G141GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n334) );
  XNOR2_X1 U373 ( .A(G22GAT), .B(G15GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n317), .B(KEYINPUT70), .ZN(n382) );
  INV_X1 U375 ( .A(n382), .ZN(n318) );
  NAND2_X1 U376 ( .A1(n318), .A2(n319), .ZN(n322) );
  INV_X1 U377 ( .A(n319), .ZN(n320) );
  NAND2_X1 U378 ( .A1(n320), .A2(n382), .ZN(n321) );
  NAND2_X1 U379 ( .A1(n322), .A2(n321), .ZN(n324) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n325), .B(KEYINPUT68), .ZN(n329) );
  XOR2_X1 U383 ( .A(G29GAT), .B(G43GAT), .Z(n327) );
  XNOR2_X1 U384 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n364) );
  XOR2_X1 U386 ( .A(n364), .B(KEYINPUT69), .Z(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U388 ( .A(G169GAT), .B(G8GAT), .Z(n408) );
  XOR2_X1 U389 ( .A(n330), .B(n408), .Z(n332) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G50GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U392 ( .A(n334), .B(n333), .Z(n453) );
  XOR2_X1 U393 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XOR2_X1 U394 ( .A(G99GAT), .B(G85GAT), .Z(n350) );
  XNOR2_X1 U395 ( .A(n436), .B(n350), .ZN(n348) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n335), .B(G148GAT), .ZN(n423) );
  NAND2_X1 U398 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n292), .B(n336), .ZN(n346) );
  XOR2_X1 U400 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n338) );
  XNOR2_X1 U401 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n383) );
  XOR2_X1 U403 ( .A(G64GAT), .B(G92GAT), .Z(n340) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n400) );
  XNOR2_X1 U406 ( .A(n383), .B(n400), .ZN(n344) );
  XOR2_X1 U407 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n342) );
  XNOR2_X1 U408 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n341) );
  XOR2_X1 U409 ( .A(n342), .B(n341), .Z(n343) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n581) );
  NAND2_X1 U411 ( .A1(n453), .A2(n552), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n349), .B(KEYINPUT46), .ZN(n387) );
  XOR2_X1 U413 ( .A(G92GAT), .B(n350), .Z(n353) );
  XNOR2_X1 U414 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n351), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U416 ( .A(G134GAT), .B(n420), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U418 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n355) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U421 ( .A(n357), .B(n356), .Z(n362) );
  XOR2_X1 U422 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n359) );
  XNOR2_X1 U423 ( .A(KEYINPUT66), .B(KEYINPUT64), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(n360), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n366) );
  XOR2_X1 U428 ( .A(G36GAT), .B(G190GAT), .Z(n365) );
  XOR2_X1 U429 ( .A(G218GAT), .B(n365), .Z(n399) );
  XNOR2_X1 U430 ( .A(n366), .B(n399), .ZN(n457) );
  INV_X1 U431 ( .A(n457), .ZN(n563) );
  XOR2_X1 U432 ( .A(G78GAT), .B(G211GAT), .Z(n368) );
  XNOR2_X1 U433 ( .A(G183GAT), .B(G127GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U435 ( .A(G64GAT), .B(G71GAT), .Z(n370) );
  XNOR2_X1 U436 ( .A(G8GAT), .B(G1GAT), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U438 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U439 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n374) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U442 ( .A(KEYINPUT77), .B(n375), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n379) );
  XNOR2_X1 U445 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U447 ( .A(n381), .B(n380), .Z(n385) );
  XNOR2_X1 U448 ( .A(n382), .B(n383), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n558) );
  XOR2_X1 U450 ( .A(G155GAT), .B(n558), .Z(n541) );
  NOR2_X1 U451 ( .A1(n563), .A2(n541), .ZN(n386) );
  AND2_X1 U452 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n388), .B(KEYINPUT47), .ZN(n395) );
  XNOR2_X1 U454 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n391) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n389), .B(n563), .ZN(n589) );
  AND2_X1 U457 ( .A1(n541), .A2(n589), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U459 ( .A1(n392), .A2(n453), .ZN(n393) );
  NAND2_X1 U460 ( .A1(n581), .A2(n393), .ZN(n394) );
  NAND2_X1 U461 ( .A1(n395), .A2(n394), .ZN(n397) );
  XNOR2_X1 U462 ( .A(KEYINPUT48), .B(KEYINPUT107), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n526) );
  XOR2_X1 U464 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U465 ( .A(G183GAT), .B(KEYINPUT18), .Z(n403) );
  XNOR2_X1 U466 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n446) );
  XNOR2_X1 U468 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n404), .B(G211GAT), .ZN(n419) );
  XNOR2_X1 U470 ( .A(n446), .B(n419), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U472 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n513), .B(KEYINPUT117), .ZN(n411) );
  NOR2_X1 U475 ( .A1(n526), .A2(n411), .ZN(n414) );
  NOR2_X1 U476 ( .A1(n529), .A2(n415), .ZN(n575) );
  XOR2_X1 U477 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n417) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U480 ( .A(n418), .B(KEYINPUT22), .Z(n422) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U483 ( .A(KEYINPUT23), .B(G218GAT), .Z(n425) );
  XNOR2_X1 U484 ( .A(G204GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U486 ( .A(n427), .B(n426), .Z(n430) );
  XNOR2_X1 U487 ( .A(G22GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n469) );
  NAND2_X1 U489 ( .A1(n575), .A2(n469), .ZN(n432) );
  INV_X1 U490 ( .A(KEYINPUT55), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n451) );
  XOR2_X1 U492 ( .A(G99GAT), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT82), .B(G176GAT), .Z(n440) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(G113GAT), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U501 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n442) );
  XNOR2_X1 U502 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U504 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n521) );
  INV_X1 U508 ( .A(n521), .ZN(n531) );
  NOR2_X1 U509 ( .A1(n451), .A2(n531), .ZN(n452) );
  XNOR2_X1 U510 ( .A(KEYINPUT119), .B(n452), .ZN(n570) );
  INV_X1 U511 ( .A(n453), .ZN(n576) );
  NOR2_X1 U512 ( .A1(n570), .A2(n576), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n454), .B(G169GAT), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(G1348GAT) );
  NOR2_X1 U516 ( .A1(n570), .A2(n457), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U518 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n469), .B(KEYINPUT67), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(KEYINPUT28), .ZN(n534) );
  XOR2_X1 U521 ( .A(n513), .B(KEYINPUT27), .Z(n527) );
  NOR2_X1 U522 ( .A1(n534), .A2(n527), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n531), .A2(n463), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n529), .A2(n464), .ZN(n476) );
  XOR2_X1 U525 ( .A(KEYINPUT95), .B(n465), .Z(n466) );
  NAND2_X1 U526 ( .A1(n469), .A2(n466), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n521), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT94), .B(n470), .Z(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT26), .B(n471), .ZN(n573) );
  NOR2_X1 U530 ( .A1(n527), .A2(n573), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n472), .A2(n529), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT96), .B(n477), .ZN(n486) );
  NOR2_X1 U535 ( .A1(n541), .A2(n486), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n589), .A2(n478), .ZN(n480) );
  NAND2_X1 U537 ( .A1(n576), .A2(n552), .ZN(n510) );
  NOR2_X1 U538 ( .A1(n497), .A2(n510), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT105), .B(n481), .Z(n523) );
  NAND2_X1 U540 ( .A1(n523), .A2(n513), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  INV_X1 U542 ( .A(n576), .ZN(n550) );
  NAND2_X1 U543 ( .A1(n550), .A2(n581), .ZN(n498) );
  INV_X1 U544 ( .A(n541), .ZN(n585) );
  NOR2_X1 U545 ( .A1(n563), .A2(n585), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U547 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT97), .B(n487), .ZN(n509) );
  NOR2_X1 U549 ( .A1(n498), .A2(n509), .ZN(n494) );
  NAND2_X1 U550 ( .A1(n529), .A2(n494), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U552 ( .A1(n494), .A2(n513), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U555 ( .A1(n494), .A2(n521), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  XOR2_X1 U558 ( .A(G22GAT), .B(KEYINPUT99), .Z(n496) );
  NAND2_X1 U559 ( .A1(n494), .A2(n534), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(KEYINPUT38), .ZN(n507) );
  NAND2_X1 U563 ( .A1(n529), .A2(n507), .ZN(n501) );
  XOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U566 ( .A1(n507), .A2(n513), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(KEYINPUT102), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n503), .ZN(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U570 ( .A1(n507), .A2(n521), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U573 ( .A1(n507), .A2(n534), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n512) );
  NOR2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n529), .A2(n516), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n516), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n534), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n529), .A2(n523), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n521), .A2(n523), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n523), .A2(n534), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT111), .Z(n537) );
  NOR2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT108), .B(n530), .ZN(n549) );
  NOR2_X1 U598 ( .A1(n531), .A2(n549), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT109), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT110), .B(n535), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n550), .A2(n544), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U605 ( .A1(n544), .A2(n552), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n544), .A2(n541), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n563), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT113), .Z(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n573), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n562), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  INV_X1 U619 ( .A(n562), .ZN(n557) );
  NOR2_X1 U620 ( .A1(n557), .A2(n567), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n557), .A2(G155GAT), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n562), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT116), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n567), .A2(n570), .ZN(n568) );
  XOR2_X1 U635 ( .A(n569), .B(n568), .Z(G1349GAT) );
  NOR2_X1 U636 ( .A1(n585), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  INV_X1 U639 ( .A(n573), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NOR2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n580) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

