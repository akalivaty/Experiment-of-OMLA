

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720;

  XNOR2_X1 U359 ( .A(n674), .B(n673), .ZN(n675) );
  INV_X1 U360 ( .A(n395), .ZN(n438) );
  INV_X1 U361 ( .A(n542), .ZN(n443) );
  NAND2_X1 U362 ( .A1(n592), .A2(n591), .ZN(n617) );
  XNOR2_X1 U363 ( .A(G101), .B(n336), .ZN(n436) );
  BUF_X1 U364 ( .A(G146), .Z(n336) );
  XNOR2_X2 U365 ( .A(n398), .B(G125), .ZN(n491) );
  XNOR2_X2 U366 ( .A(KEYINPUT76), .B(KEYINPUT33), .ZN(n348) );
  XOR2_X2 U367 ( .A(n663), .B(n662), .Z(n351) );
  INV_X2 U368 ( .A(KEYINPUT86), .ZN(n453) );
  XNOR2_X2 U369 ( .A(n541), .B(n348), .ZN(n395) );
  XOR2_X1 U370 ( .A(n523), .B(n522), .Z(n337) );
  AND2_X2 U371 ( .A1(n365), .A2(n363), .ZN(n362) );
  INV_X2 U372 ( .A(KEYINPUT4), .ZN(n425) );
  NAND2_X2 U373 ( .A1(n455), .A2(n454), .ZN(n457) );
  OR2_X2 U374 ( .A1(n476), .A2(G902), .ZN(n477) );
  NOR2_X2 U375 ( .A1(n590), .A2(n502), .ZN(n420) );
  NOR2_X2 U376 ( .A1(n661), .A2(n603), .ZN(n499) );
  AND2_X1 U377 ( .A1(n361), .A2(n360), .ZN(n359) );
  NOR2_X2 U378 ( .A1(n714), .A2(n720), .ZN(n422) );
  INV_X1 U379 ( .A(n583), .ZN(n554) );
  AND2_X1 U380 ( .A1(n444), .A2(n440), .ZN(n439) );
  NOR2_X1 U381 ( .A1(n438), .A2(n394), .ZN(n660) );
  XNOR2_X1 U382 ( .A(n420), .B(n421), .ZN(n547) );
  AND2_X1 U383 ( .A1(n648), .A2(n585), .ZN(n578) );
  XNOR2_X1 U384 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U385 ( .A(n390), .B(n399), .ZN(n497) );
  XNOR2_X1 U386 ( .A(n415), .B(n494), .ZN(n695) );
  XNOR2_X2 U387 ( .A(G104), .B(G110), .ZN(n449) );
  INV_X2 U388 ( .A(G953), .ZN(n709) );
  INV_X1 U389 ( .A(G146), .ZN(n398) );
  NAND2_X2 U390 ( .A1(n567), .A2(n633), .ZN(n586) );
  AND2_X2 U391 ( .A1(n427), .A2(n426), .ZN(n602) );
  XNOR2_X1 U392 ( .A(n560), .B(n349), .ZN(n355) );
  NAND2_X1 U393 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U394 ( .A1(n579), .A2(n646), .ZN(n566) );
  XNOR2_X1 U395 ( .A(n449), .B(G107), .ZN(n493) );
  XNOR2_X1 U396 ( .A(G131), .B(KEYINPUT73), .ZN(n520) );
  XNOR2_X1 U397 ( .A(n378), .B(n377), .ZN(n494) );
  XNOR2_X1 U398 ( .A(G116), .B(KEYINPUT3), .ZN(n377) );
  XNOR2_X1 U399 ( .A(n448), .B(G119), .ZN(n378) );
  INV_X1 U400 ( .A(G113), .ZN(n448) );
  XNOR2_X1 U401 ( .A(n491), .B(n410), .ZN(n518) );
  INV_X1 U402 ( .A(KEYINPUT10), .ZN(n410) );
  XNOR2_X1 U403 ( .A(n385), .B(KEYINPUT50), .ZN(n384) );
  INV_X1 U404 ( .A(KEYINPUT115), .ZN(n385) );
  XNOR2_X1 U405 ( .A(G140), .B(KEYINPUT97), .ZN(n522) );
  XOR2_X1 U406 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n523) );
  XNOR2_X1 U407 ( .A(n459), .B(G137), .ZN(n376) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(KEYINPUT5), .Z(n459) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n517) );
  XOR2_X1 U410 ( .A(KEYINPUT7), .B(G107), .Z(n504) );
  XNOR2_X1 U411 ( .A(G116), .B(G122), .ZN(n503) );
  XOR2_X1 U412 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n506) );
  XOR2_X1 U413 ( .A(G137), .B(G140), .Z(n479) );
  XNOR2_X1 U414 ( .A(n347), .B(n496), .ZN(n399) );
  XNOR2_X1 U415 ( .A(n495), .B(G101), .ZN(n496) );
  INV_X1 U416 ( .A(KEYINPUT81), .ZN(n495) );
  XOR2_X1 U417 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n492) );
  XNOR2_X1 U418 ( .A(n423), .B(KEYINPUT105), .ZN(n631) );
  INV_X1 U419 ( .A(KEYINPUT30), .ZN(n409) );
  INV_X1 U420 ( .A(n478), .ZN(n648) );
  XNOR2_X1 U421 ( .A(n493), .B(n345), .ZN(n415) );
  XNOR2_X1 U422 ( .A(KEYINPUT93), .B(KEYINPUT75), .ZN(n467) );
  XNOR2_X1 U423 ( .A(G119), .B(G128), .ZN(n465) );
  XNOR2_X1 U424 ( .A(n434), .B(n433), .ZN(n509) );
  INV_X1 U425 ( .A(KEYINPUT8), .ZN(n433) );
  NAND2_X1 U426 ( .A1(n709), .A2(G234), .ZN(n434) );
  XOR2_X1 U427 ( .A(n528), .B(n527), .Z(n674) );
  XNOR2_X1 U428 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U429 ( .A(G113), .B(G143), .ZN(n515) );
  XNOR2_X1 U430 ( .A(n569), .B(n568), .ZN(n573) );
  INV_X1 U431 ( .A(n543), .ZN(n442) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n372) );
  INV_X1 U433 ( .A(KEYINPUT84), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n432), .B(n431), .ZN(n539) );
  XNOR2_X1 U435 ( .A(n475), .B(KEYINPUT25), .ZN(n431) );
  NOR2_X1 U436 ( .A1(n683), .A2(G902), .ZN(n432) );
  XNOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT22), .ZN(n534) );
  NOR2_X1 U438 ( .A1(G952), .A2(n709), .ZN(n688) );
  XNOR2_X1 U439 ( .A(n369), .B(KEYINPUT47), .ZN(n407) );
  INV_X2 U440 ( .A(G128), .ZN(n452) );
  NOR2_X1 U441 ( .A1(n472), .A2(KEYINPUT88), .ZN(n364) );
  NAND2_X1 U442 ( .A1(n386), .A2(n383), .ZN(n650) );
  AND2_X1 U443 ( .A1(n649), .A2(n478), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n647), .B(n384), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n371), .B(KEYINPUT44), .ZN(n559) );
  XNOR2_X1 U446 ( .A(n524), .B(n337), .ZN(n525) );
  XNOR2_X1 U447 ( .A(n518), .B(n519), .ZN(n526) );
  XOR2_X1 U448 ( .A(G104), .B(G122), .Z(n516) );
  NAND2_X1 U449 ( .A1(n472), .A2(KEYINPUT88), .ZN(n360) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n486) );
  OR2_X1 U451 ( .A1(G237), .A2(G902), .ZN(n500) );
  INV_X1 U452 ( .A(KEYINPUT38), .ZN(n424) );
  NOR2_X1 U453 ( .A1(n577), .A2(n576), .ZN(n585) );
  XNOR2_X1 U454 ( .A(n446), .B(n540), .ZN(n358) );
  INV_X1 U455 ( .A(KEYINPUT79), .ZN(n540) );
  NOR2_X1 U456 ( .A1(n645), .A2(n646), .ZN(n446) );
  XNOR2_X1 U457 ( .A(n579), .B(n447), .ZN(n645) );
  XNOR2_X1 U458 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n447) );
  INV_X1 U459 ( .A(KEYINPUT0), .ZN(n421) );
  XNOR2_X1 U460 ( .A(n483), .B(n462), .ZN(n476) );
  XNOR2_X1 U461 ( .A(n494), .B(n376), .ZN(n461) );
  INV_X1 U462 ( .A(n713), .ZN(n426) );
  INV_X1 U463 ( .A(G134), .ZN(n458) );
  XNOR2_X1 U464 ( .A(KEYINPUT99), .B(KEYINPUT101), .ZN(n505) );
  XNOR2_X1 U465 ( .A(n416), .B(n695), .ZN(n661) );
  XNOR2_X1 U466 ( .A(n396), .B(n497), .ZN(n416) );
  AND2_X1 U467 ( .A1(n379), .A2(n340), .ZN(n654) );
  XNOR2_X1 U468 ( .A(n380), .B(KEYINPUT116), .ZN(n379) );
  AND2_X1 U469 ( .A1(n441), .A2(n544), .ZN(n440) );
  AND2_X1 U470 ( .A1(n566), .A2(n401), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n565), .B(n409), .ZN(n408) );
  INV_X1 U472 ( .A(n577), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n530), .B(n529), .ZN(n551) );
  XNOR2_X1 U474 ( .A(KEYINPUT13), .B(G475), .ZN(n529) );
  XNOR2_X1 U475 ( .A(n471), .B(n700), .ZN(n683) );
  XNOR2_X1 U476 ( .A(n370), .B(n346), .ZN(n471) );
  XNOR2_X1 U477 ( .A(n470), .B(n469), .ZN(n370) );
  INV_X1 U478 ( .A(n653), .ZN(n394) );
  XNOR2_X1 U479 ( .A(n581), .B(n582), .ZN(n714) );
  XNOR2_X1 U480 ( .A(n538), .B(KEYINPUT67), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n338), .A2(n392), .ZN(n391) );
  NAND2_X1 U482 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U483 ( .A(n688), .ZN(n412) );
  XNOR2_X1 U484 ( .A(n414), .B(n350), .ZN(n413) );
  XNOR2_X1 U485 ( .A(n388), .B(n387), .ZN(G75) );
  XNOR2_X1 U486 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n387) );
  NAND2_X1 U487 ( .A1(n339), .A2(n389), .ZN(n388) );
  NOR2_X1 U488 ( .A1(n660), .A2(G953), .ZN(n389) );
  OR2_X1 U489 ( .A1(n402), .A2(n539), .ZN(n338) );
  AND2_X1 U490 ( .A1(n659), .A2(n658), .ZN(n339) );
  XOR2_X1 U491 ( .A(KEYINPUT119), .B(n641), .Z(n340) );
  AND2_X1 U492 ( .A1(n408), .A2(n400), .ZN(n341) );
  XOR2_X1 U493 ( .A(KEYINPUT87), .B(n616), .Z(n342) );
  XNOR2_X1 U494 ( .A(n575), .B(KEYINPUT103), .ZN(n343) );
  BUF_X1 U495 ( .A(n645), .Z(n405) );
  AND2_X1 U496 ( .A1(n542), .A2(n543), .ZN(n344) );
  XOR2_X1 U497 ( .A(G122), .B(KEYINPUT16), .Z(n345) );
  AND2_X1 U498 ( .A1(G221), .A2(n509), .ZN(n346) );
  AND2_X1 U499 ( .A1(G224), .A2(n709), .ZN(n347) );
  BUF_X1 U500 ( .A(n648), .Z(n402) );
  NOR2_X1 U501 ( .A1(n549), .A2(n551), .ZN(n580) );
  XOR2_X1 U502 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n349) );
  XOR2_X1 U503 ( .A(n464), .B(n463), .Z(n350) );
  XOR2_X1 U504 ( .A(KEYINPUT15), .B(G902), .Z(n603) );
  XOR2_X1 U505 ( .A(n596), .B(KEYINPUT48), .Z(n352) );
  NAND2_X1 U506 ( .A1(n438), .A2(n442), .ZN(n437) );
  OR2_X2 U507 ( .A1(n547), .A2(n451), .ZN(n450) );
  BUF_X1 U508 ( .A(n358), .Z(n353) );
  NAND2_X1 U509 ( .A1(n634), .A2(n633), .ZN(n423) );
  XNOR2_X1 U510 ( .A(n445), .B(KEYINPUT35), .ZN(n715) );
  NAND2_X1 U511 ( .A1(n439), .A2(n437), .ZN(n445) );
  NAND2_X1 U512 ( .A1(n358), .A2(n554), .ZN(n541) );
  NAND2_X1 U513 ( .A1(n537), .A2(n372), .ZN(n418) );
  XNOR2_X1 U514 ( .A(n567), .B(n424), .ZN(n634) );
  INV_X1 U515 ( .A(n438), .ZN(n354) );
  BUF_X1 U516 ( .A(n579), .Z(n356) );
  XNOR2_X1 U517 ( .A(n560), .B(n349), .ZN(n692) );
  BUF_X1 U518 ( .A(n672), .Z(n684) );
  NAND2_X1 U519 ( .A1(n672), .A2(G472), .ZN(n414) );
  BUF_X1 U520 ( .A(n513), .Z(n357) );
  NAND2_X1 U521 ( .A1(n353), .A2(n402), .ZN(n651) );
  NOR2_X1 U522 ( .A1(n355), .A2(n707), .ZN(n604) );
  NAND2_X1 U523 ( .A1(n362), .A2(n359), .ZN(n605) );
  NAND2_X1 U524 ( .A1(n707), .A2(n364), .ZN(n361) );
  NAND2_X1 U525 ( .A1(n692), .A2(n364), .ZN(n363) );
  NAND2_X1 U526 ( .A1(n366), .A2(n367), .ZN(n365) );
  INV_X1 U527 ( .A(n355), .ZN(n366) );
  NOR2_X1 U528 ( .A1(n707), .A2(n603), .ZN(n367) );
  NAND2_X2 U529 ( .A1(n602), .A2(n629), .ZN(n707) );
  XNOR2_X1 U530 ( .A(n491), .B(n492), .ZN(n397) );
  XNOR2_X2 U531 ( .A(n368), .B(KEYINPUT41), .ZN(n653) );
  NAND2_X1 U532 ( .A1(n631), .A2(n580), .ZN(n368) );
  NOR2_X1 U533 ( .A1(n573), .A2(n620), .ZN(n574) );
  NAND2_X1 U534 ( .A1(n594), .A2(KEYINPUT72), .ZN(n369) );
  NOR2_X2 U535 ( .A1(n715), .A2(n545), .ZN(n371) );
  NAND2_X1 U536 ( .A1(n537), .A2(n405), .ZN(n553) );
  NAND2_X1 U537 ( .A1(n536), .A2(n375), .ZN(n374) );
  NOR2_X1 U538 ( .A1(n405), .A2(n343), .ZN(n375) );
  NAND2_X1 U539 ( .A1(n381), .A2(n653), .ZN(n380) );
  XNOR2_X1 U540 ( .A(n652), .B(n382), .ZN(n381) );
  INV_X1 U541 ( .A(KEYINPUT51), .ZN(n382) );
  XNOR2_X1 U542 ( .A(n390), .B(n436), .ZN(n435) );
  XNOR2_X2 U543 ( .A(n702), .B(KEYINPUT71), .ZN(n390) );
  NAND2_X1 U544 ( .A1(n537), .A2(n391), .ZN(n419) );
  INV_X1 U545 ( .A(n405), .ZN(n392) );
  XNOR2_X2 U546 ( .A(n450), .B(n534), .ZN(n537) );
  XNOR2_X1 U547 ( .A(n393), .B(n397), .ZN(n396) );
  XNOR2_X2 U548 ( .A(n393), .B(n458), .ZN(n513) );
  XNOR2_X2 U549 ( .A(n457), .B(n456), .ZN(n393) );
  NAND2_X1 U550 ( .A1(n395), .A2(n344), .ZN(n444) );
  NAND2_X1 U551 ( .A1(n640), .A2(n354), .ZN(n641) );
  XNOR2_X2 U552 ( .A(n586), .B(n501), .ZN(n590) );
  XNOR2_X1 U553 ( .A(n554), .B(KEYINPUT85), .ZN(n536) );
  NOR2_X2 U554 ( .A1(n617), .A2(n593), .ZN(n594) );
  AND2_X2 U555 ( .A1(n404), .A2(n403), .ZN(n592) );
  INV_X1 U556 ( .A(n356), .ZN(n403) );
  XNOR2_X1 U557 ( .A(n578), .B(KEYINPUT28), .ZN(n404) );
  XNOR2_X1 U558 ( .A(n422), .B(KEYINPUT46), .ZN(n430) );
  NAND2_X1 U559 ( .A1(n672), .A2(G210), .ZN(n664) );
  XNOR2_X2 U560 ( .A(n606), .B(KEYINPUT66), .ZN(n672) );
  XNOR2_X1 U561 ( .A(n406), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U562 ( .A1(n665), .A2(n688), .ZN(n406) );
  NOR2_X1 U563 ( .A1(n407), .A2(n626), .ZN(n595) );
  XNOR2_X1 U564 ( .A(n428), .B(n352), .ZN(n427) );
  XNOR2_X1 U565 ( .A(n411), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U566 ( .A1(n672), .A2(G475), .ZN(n676) );
  NOR2_X2 U567 ( .A1(n677), .A2(n688), .ZN(n679) );
  NAND2_X1 U568 ( .A1(n580), .A2(n642), .ZN(n451) );
  NAND2_X1 U569 ( .A1(n719), .A2(n717), .ZN(n545) );
  XNOR2_X2 U570 ( .A(n418), .B(n417), .ZN(n717) );
  XNOR2_X2 U571 ( .A(n419), .B(KEYINPUT104), .ZN(n719) );
  INV_X1 U572 ( .A(n567), .ZN(n600) );
  XNOR2_X2 U573 ( .A(n425), .B(KEYINPUT65), .ZN(n702) );
  NAND2_X1 U574 ( .A1(n430), .A2(n429), .ZN(n428) );
  AND2_X1 U575 ( .A1(n595), .A2(n342), .ZN(n429) );
  XNOR2_X2 U576 ( .A(n701), .B(n435), .ZN(n483) );
  XNOR2_X2 U577 ( .A(n513), .B(n520), .ZN(n701) );
  NAND2_X1 U578 ( .A1(n443), .A2(n442), .ZN(n441) );
  XNOR2_X1 U579 ( .A(n664), .B(n351), .ZN(n665) );
  XNOR2_X2 U580 ( .A(n499), .B(n498), .ZN(n567) );
  INV_X1 U581 ( .A(KEYINPUT89), .ZN(n596) );
  XNOR2_X1 U582 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U583 ( .A(G143), .ZN(n456) );
  XNOR2_X1 U584 ( .A(G469), .B(KEYINPUT74), .ZN(n484) );
  INV_X1 U585 ( .A(KEYINPUT39), .ZN(n568) );
  XNOR2_X1 U586 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U587 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(KEYINPUT62), .Z(n464) );
  NAND2_X1 U589 ( .A1(n452), .A2(KEYINPUT86), .ZN(n455) );
  NAND2_X1 U590 ( .A1(n453), .A2(G128), .ZN(n454) );
  AND2_X1 U591 ( .A1(n517), .A2(G210), .ZN(n460) );
  XNOR2_X1 U592 ( .A(n476), .B(KEYINPUT109), .ZN(n463) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(G110), .Z(n466) );
  XNOR2_X1 U594 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U595 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n468) );
  XNOR2_X1 U596 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U597 ( .A(n479), .B(n518), .ZN(n700) );
  XOR2_X1 U598 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n474) );
  INV_X1 U599 ( .A(n603), .ZN(n472) );
  NAND2_X1 U600 ( .A1(G234), .A2(n472), .ZN(n473) );
  XNOR2_X1 U601 ( .A(n474), .B(n473), .ZN(n531) );
  NAND2_X1 U602 ( .A1(G217), .A2(n531), .ZN(n475) );
  INV_X1 U603 ( .A(n539), .ZN(n575) );
  XNOR2_X2 U604 ( .A(n477), .B(G472), .ZN(n564) );
  INV_X1 U605 ( .A(n564), .ZN(n478) );
  XOR2_X1 U606 ( .A(n493), .B(n479), .Z(n481) );
  NAND2_X1 U607 ( .A1(G227), .A2(n709), .ZN(n480) );
  XNOR2_X1 U608 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U609 ( .A(n483), .B(n482), .ZN(n666) );
  NOR2_X1 U610 ( .A1(n666), .A2(G902), .ZN(n485) );
  XNOR2_X2 U611 ( .A(n485), .B(n484), .ZN(n579) );
  XNOR2_X1 U612 ( .A(n486), .B(KEYINPUT14), .ZN(n487) );
  XNOR2_X1 U613 ( .A(KEYINPUT78), .B(n487), .ZN(n488) );
  NAND2_X1 U614 ( .A1(G952), .A2(n488), .ZN(n656) );
  NOR2_X1 U615 ( .A1(G953), .A2(n656), .ZN(n563) );
  AND2_X1 U616 ( .A1(n488), .A2(G953), .ZN(n489) );
  NAND2_X1 U617 ( .A1(G902), .A2(n489), .ZN(n561) );
  NOR2_X1 U618 ( .A1(G898), .A2(n561), .ZN(n490) );
  NOR2_X1 U619 ( .A1(n563), .A2(n490), .ZN(n502) );
  XNOR2_X1 U620 ( .A(KEYINPUT19), .B(KEYINPUT69), .ZN(n501) );
  NAND2_X1 U621 ( .A1(G210), .A2(n500), .ZN(n498) );
  NAND2_X1 U622 ( .A1(G214), .A2(n500), .ZN(n633) );
  XNOR2_X1 U623 ( .A(n504), .B(n503), .ZN(n508) );
  XNOR2_X1 U624 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U625 ( .A(n508), .B(n507), .Z(n511) );
  NAND2_X1 U626 ( .A1(G217), .A2(n509), .ZN(n510) );
  XNOR2_X1 U627 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U628 ( .A(n357), .B(n512), .ZN(n681) );
  NOR2_X1 U629 ( .A1(G902), .A2(n681), .ZN(n514) );
  XOR2_X1 U630 ( .A(G478), .B(n514), .Z(n549) );
  XNOR2_X1 U631 ( .A(n516), .B(n515), .ZN(n528) );
  NAND2_X1 U632 ( .A1(G214), .A2(n517), .ZN(n519) );
  INV_X1 U633 ( .A(n520), .ZN(n521) );
  XNOR2_X1 U634 ( .A(n521), .B(KEYINPUT98), .ZN(n524) );
  NOR2_X1 U635 ( .A1(G902), .A2(n674), .ZN(n530) );
  INV_X1 U636 ( .A(n580), .ZN(n636) );
  XOR2_X1 U637 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n533) );
  NAND2_X1 U638 ( .A1(n531), .A2(G221), .ZN(n532) );
  XNOR2_X1 U639 ( .A(n533), .B(n532), .ZN(n642) );
  XNOR2_X1 U640 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n535) );
  XNOR2_X1 U641 ( .A(n535), .B(n564), .ZN(n583) );
  XNOR2_X1 U642 ( .A(KEYINPUT83), .B(KEYINPUT32), .ZN(n538) );
  INV_X1 U643 ( .A(n547), .ZN(n542) );
  NAND2_X1 U644 ( .A1(n642), .A2(n539), .ZN(n646) );
  XOR2_X1 U645 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n543) );
  NAND2_X1 U646 ( .A1(n549), .A2(n551), .ZN(n571) );
  INV_X1 U647 ( .A(n571), .ZN(n544) );
  NOR2_X1 U648 ( .A1(n402), .A2(n443), .ZN(n546) );
  NAND2_X1 U649 ( .A1(n566), .A2(n546), .ZN(n611) );
  NOR2_X1 U650 ( .A1(n443), .A2(n651), .ZN(n548) );
  XNOR2_X1 U651 ( .A(n548), .B(KEYINPUT31), .ZN(n622) );
  NAND2_X1 U652 ( .A1(n611), .A2(n622), .ZN(n552) );
  INV_X1 U653 ( .A(n549), .ZN(n550) );
  OR2_X1 U654 ( .A1(n550), .A2(n551), .ZN(n623) );
  NAND2_X1 U655 ( .A1(n551), .A2(n550), .ZN(n620) );
  NAND2_X1 U656 ( .A1(n623), .A2(n620), .ZN(n630) );
  NAND2_X1 U657 ( .A1(n552), .A2(n630), .ZN(n557) );
  NOR2_X1 U658 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U659 ( .A(n555), .B(KEYINPUT90), .ZN(n556) );
  NAND2_X1 U660 ( .A1(n556), .A2(n343), .ZN(n607) );
  AND2_X1 U661 ( .A1(n557), .A2(n607), .ZN(n558) );
  NOR2_X1 U662 ( .A1(G900), .A2(n561), .ZN(n562) );
  NOR2_X1 U663 ( .A1(n563), .A2(n562), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n564), .A2(n633), .ZN(n565) );
  NAND2_X1 U665 ( .A1(n341), .A2(n634), .ZN(n569) );
  OR2_X1 U666 ( .A1(n573), .A2(n623), .ZN(n570) );
  XNOR2_X1 U667 ( .A(n570), .B(KEYINPUT107), .ZN(n713) );
  NOR2_X1 U668 ( .A1(n600), .A2(n571), .ZN(n572) );
  NAND2_X1 U669 ( .A1(n341), .A2(n572), .ZN(n616) );
  XNOR2_X1 U670 ( .A(n574), .B(KEYINPUT40), .ZN(n720) );
  XOR2_X1 U671 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n582) );
  NAND2_X1 U672 ( .A1(n642), .A2(n575), .ZN(n576) );
  NAND2_X1 U673 ( .A1(n592), .A2(n653), .ZN(n581) );
  NOR2_X1 U674 ( .A1(n583), .A2(n620), .ZN(n584) );
  NAND2_X1 U675 ( .A1(n585), .A2(n584), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n586), .A2(n597), .ZN(n588) );
  XNOR2_X1 U677 ( .A(KEYINPUT36), .B(KEYINPUT91), .ZN(n587) );
  XNOR2_X1 U678 ( .A(n588), .B(n587), .ZN(n589) );
  NOR2_X1 U679 ( .A1(n405), .A2(n589), .ZN(n626) );
  INV_X1 U680 ( .A(n590), .ZN(n591) );
  INV_X1 U681 ( .A(n630), .ZN(n593) );
  NOR2_X1 U682 ( .A1(n392), .A2(n597), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n598), .A2(n633), .ZN(n599) );
  XNOR2_X1 U684 ( .A(n599), .B(KEYINPUT43), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n629) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT2), .ZN(n659) );
  NOR2_X2 U687 ( .A1(n605), .A2(n659), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n607), .B(G101), .ZN(G3) );
  NOR2_X1 U689 ( .A1(n620), .A2(n611), .ZN(n608) );
  XOR2_X1 U690 ( .A(G104), .B(n608), .Z(G6) );
  XOR2_X1 U691 ( .A(KEYINPUT26), .B(KEYINPUT110), .Z(n610) );
  XNOR2_X1 U692 ( .A(G107), .B(KEYINPUT27), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n610), .B(n609), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n623), .A2(n611), .ZN(n612) );
  XOR2_X1 U695 ( .A(n613), .B(n612), .Z(G9) );
  NOR2_X1 U696 ( .A1(n623), .A2(n617), .ZN(n615) );
  XNOR2_X1 U697 ( .A(G128), .B(KEYINPUT29), .ZN(n614) );
  XNOR2_X1 U698 ( .A(n615), .B(n614), .ZN(G30) );
  XNOR2_X1 U699 ( .A(G143), .B(n616), .ZN(G45) );
  NOR2_X1 U700 ( .A1(n620), .A2(n617), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n336), .B(KEYINPUT111), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n619), .B(n618), .ZN(G48) );
  NOR2_X1 U703 ( .A1(n620), .A2(n622), .ZN(n621) );
  XOR2_X1 U704 ( .A(G113), .B(n621), .Z(G15) );
  NOR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U706 ( .A(KEYINPUT112), .B(n624), .Z(n625) );
  XNOR2_X1 U707 ( .A(G116), .B(n625), .ZN(G18) );
  XOR2_X1 U708 ( .A(KEYINPUT113), .B(KEYINPUT37), .Z(n628) );
  XNOR2_X1 U709 ( .A(G125), .B(n626), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n628), .B(n627), .ZN(G27) );
  XNOR2_X1 U711 ( .A(G140), .B(n629), .ZN(G42) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U713 ( .A(KEYINPUT117), .B(n632), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U717 ( .A(KEYINPUT118), .B(n639), .Z(n640) );
  NOR2_X1 U718 ( .A1(n642), .A2(n343), .ZN(n644) );
  XNOR2_X1 U719 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n644), .B(n643), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n646), .A2(n405), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT52), .B(n654), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT120), .B(n657), .Z(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n663) );
  XNOR2_X1 U727 ( .A(n661), .B(KEYINPUT92), .ZN(n662) );
  NAND2_X1 U728 ( .A1(G469), .A2(n684), .ZN(n670) );
  BUF_X1 U729 ( .A(n666), .Z(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n667) );
  NOR2_X1 U731 ( .A1(n688), .A2(n671), .ZN(G54) );
  XOR2_X1 U732 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n673) );
  XNOR2_X1 U733 ( .A(KEYINPUT70), .B(KEYINPUT60), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n679), .B(n678), .ZN(G60) );
  NAND2_X1 U735 ( .A1(G478), .A2(n684), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U737 ( .A1(n682), .A2(n688), .ZN(G63) );
  XOR2_X1 U738 ( .A(n683), .B(KEYINPUT123), .Z(n686) );
  NAND2_X1 U739 ( .A1(G217), .A2(n684), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U741 ( .A1(n687), .A2(n688), .ZN(G66) );
  NAND2_X1 U742 ( .A1(G953), .A2(G224), .ZN(n689) );
  XNOR2_X1 U743 ( .A(KEYINPUT61), .B(n689), .ZN(n690) );
  NAND2_X1 U744 ( .A1(n690), .A2(G898), .ZN(n691) );
  XOR2_X1 U745 ( .A(KEYINPUT124), .B(n691), .Z(n694) );
  NOR2_X1 U746 ( .A1(G953), .A2(n692), .ZN(n693) );
  NOR2_X1 U747 ( .A1(n694), .A2(n693), .ZN(n699) );
  XNOR2_X1 U748 ( .A(n695), .B(G101), .ZN(n697) );
  NOR2_X1 U749 ( .A1(n709), .A2(G898), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U751 ( .A(n699), .B(n698), .Z(G69) );
  XNOR2_X1 U752 ( .A(n700), .B(KEYINPUT125), .ZN(n704) );
  XNOR2_X1 U753 ( .A(n701), .B(n702), .ZN(n703) );
  XOR2_X1 U754 ( .A(n704), .B(n703), .Z(n708) );
  XNOR2_X1 U755 ( .A(G227), .B(n708), .ZN(n705) );
  NAND2_X1 U756 ( .A1(G900), .A2(n705), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n706), .A2(G953), .ZN(n712) );
  XNOR2_X1 U758 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U759 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U760 ( .A1(n712), .A2(n711), .ZN(G72) );
  XOR2_X1 U761 ( .A(G134), .B(n713), .Z(G36) );
  XOR2_X1 U762 ( .A(n714), .B(G137), .Z(G39) );
  BUF_X1 U763 ( .A(n715), .Z(n716) );
  XOR2_X1 U764 ( .A(G122), .B(n716), .Z(G24) );
  XNOR2_X1 U765 ( .A(n717), .B(G119), .ZN(n718) );
  XNOR2_X1 U766 ( .A(n718), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U767 ( .A(n719), .B(G110), .ZN(G12) );
  XOR2_X1 U768 ( .A(n720), .B(G131), .Z(G33) );
endmodule

