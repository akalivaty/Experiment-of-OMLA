//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT93), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G122), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT69), .B1(new_n194), .B2(G116), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n192), .A3(G119), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT2), .B(G113), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(KEYINPUT70), .A3(new_n200), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT70), .B1(new_n198), .B2(new_n200), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(G101), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n208), .A2(new_n211), .A3(new_n217), .A4(new_n212), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n206), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n221));
  INV_X1    g035(.A(new_n193), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n196), .B1(new_n192), .B2(G119), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n194), .A2(KEYINPUT69), .A3(G116), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n225), .B2(new_n199), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n203), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n228), .A2(KEYINPUT5), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(KEYINPUT5), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT90), .B1(new_n231), .B2(new_n222), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n198), .A2(new_n231), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n234), .A3(new_n193), .A4(new_n230), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(new_n233), .A3(G113), .A4(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n207), .A2(G107), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n210), .A2(G104), .ZN(new_n238));
  OAI21_X1  g052(.A(G101), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT85), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT85), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n218), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n227), .A2(new_n236), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n191), .B1(new_n220), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT6), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT91), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n220), .A2(new_n244), .A3(new_n191), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT6), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n247), .B(new_n248), .C1(new_n250), .C2(new_n245), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n220), .A2(new_n244), .ZN(new_n252));
  INV_X1    g066(.A(new_n191), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n254), .A2(new_n249), .A3(KEYINPUT91), .A4(KEYINPUT6), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n257), .B2(G146), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(G146), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  OAI211_X1 g075(.A(G128), .B(new_n258), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(G146), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n263), .B(new_n264), .C1(KEYINPUT1), .C2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT0), .A3(G128), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G224), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n256), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n276), .A2(KEYINPUT7), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT92), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n280), .A2(KEYINPUT92), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n274), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n249), .B(new_n283), .C1(new_n285), .C2(new_n282), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n191), .B(KEYINPUT8), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n227), .A2(new_n236), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n240), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n291), .A2(G113), .A3(new_n232), .A4(new_n235), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n292), .A2(new_n227), .A3(new_n218), .A4(new_n239), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n288), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n279), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n190), .B1(new_n278), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n277), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n251), .B2(new_n255), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n299), .A2(new_n189), .A3(new_n295), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n187), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT94), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n278), .A2(new_n190), .A3(new_n296), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n189), .B1(new_n299), .B2(new_n295), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n187), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT100), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G122), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT14), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(KEYINPUT98), .A3(G107), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT98), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n192), .A2(G122), .ZN(new_n315));
  INV_X1    g129(.A(G122), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n315), .A2(new_n317), .A3(new_n310), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n312), .A2(G107), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT96), .B1(new_n257), .B2(G128), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT96), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n265), .A3(G143), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n257), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G134), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n329), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n309), .A2(new_n210), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n321), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT99), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT99), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n321), .A2(new_n331), .A3(new_n335), .A4(new_n332), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT13), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n322), .A2(new_n324), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT97), .ZN(new_n339));
  OAI22_X1  g153(.A1(new_n338), .A2(new_n339), .B1(new_n337), .B2(new_n326), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n338), .A2(new_n339), .ZN(new_n341));
  OAI21_X1  g155(.A(G134), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n309), .B(new_n210), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(new_n330), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n336), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT9), .B(G234), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT78), .B(G217), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n275), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n333), .A2(KEYINPUT99), .B1(new_n342), .B2(new_n344), .ZN(new_n352));
  INV_X1    g166(.A(new_n350), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n336), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT75), .B(G902), .ZN(new_n356));
  INV_X1    g170(.A(G478), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT15), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n355), .B2(new_n356), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n308), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n360), .A3(KEYINPUT100), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G952), .ZN(new_n367));
  AOI211_X1 g181(.A(G953), .B(new_n367), .C1(G234), .C2(G237), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n275), .B(new_n356), .C1(G234), .C2(G237), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT21), .B(G898), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n275), .A3(G214), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(G143), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT18), .ZN(new_n375));
  INV_X1    g189(.A(G131), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n373), .B(new_n257), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT18), .A3(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(G125), .B(G140), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n260), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(G131), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n374), .A2(new_n376), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(KEYINPUT17), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n268), .A2(KEYINPUT16), .A3(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n260), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(G146), .A3(new_n388), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(new_n391), .C1(new_n383), .C2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n382), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G113), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n207), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n394), .B(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G475), .B1(new_n397), .B2(G902), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n396), .B(new_n382), .C1(new_n386), .C2(new_n393), .ZN(new_n399));
  INV_X1    g213(.A(new_n382), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n380), .A2(KEYINPUT19), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n380), .A2(KEYINPUT19), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n260), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n387), .A2(new_n405), .A3(G146), .A4(new_n388), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n407), .A2(KEYINPUT95), .B1(new_n383), .B2(new_n384), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT95), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n401), .A2(new_n404), .A3(new_n409), .A4(new_n406), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n400), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n399), .B1(new_n411), .B2(new_n396), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n398), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n366), .A2(new_n371), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n302), .A2(new_n307), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n279), .ZN(new_n422));
  INV_X1    g236(.A(new_n356), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT11), .B1(new_n329), .B2(G137), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT11), .ZN(new_n425));
  INV_X1    g239(.A(G137), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G134), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n426), .B2(G134), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n329), .A2(KEYINPUT65), .A3(G137), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G131), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n424), .A2(new_n427), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n435), .A2(new_n376), .A3(new_n430), .A4(new_n431), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT66), .B(G131), .C1(new_n428), .C2(new_n432), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n262), .A2(new_n266), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n240), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n262), .A2(new_n218), .A3(new_n239), .A4(new_n266), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(KEYINPUT12), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT12), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n437), .A2(new_n438), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n441), .A2(new_n442), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n448), .A3(KEYINPUT88), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n446), .A2(KEYINPUT86), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n437), .B2(new_n438), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n273), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n219), .A3(new_n215), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n241), .A2(new_n267), .A3(KEYINPUT10), .A4(new_n243), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT10), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n442), .A2(KEYINPUT84), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT84), .B1(new_n442), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n458), .B(new_n459), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  INV_X1    g280(.A(G227), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G953), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n466), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n451), .A2(new_n452), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n463), .A2(new_n453), .A3(new_n455), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n463), .A2(new_n439), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n469), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n423), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n422), .B1(new_n476), .B2(new_n421), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n465), .A2(new_n470), .A3(new_n473), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n470), .B1(new_n465), .B2(new_n449), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT87), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n472), .B1(new_n444), .B2(new_n448), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(new_n478), .C1(new_n483), .C2(new_n470), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n484), .A3(G469), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G221), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n348), .B2(new_n279), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n488), .B(KEYINPUT83), .Z(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n420), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n329), .B2(G137), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n329), .A2(G137), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n426), .A2(KEYINPUT67), .A3(G134), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n436), .A2(new_n499), .A3(new_n266), .A4(new_n262), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n267), .A2(KEYINPUT68), .A3(new_n436), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n437), .A2(new_n438), .A3(new_n457), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n206), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n206), .A2(KEYINPUT72), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n201), .B1(new_n226), .B2(new_n203), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n508), .A2(new_n511), .A3(new_n505), .A4(new_n500), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n493), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n512), .A2(new_n493), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n372), .A2(new_n275), .A3(G210), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT27), .Z(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT26), .B(G101), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n517), .B(new_n518), .Z(new_n519));
  NOR2_X1   g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n512), .A2(new_n519), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n506), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n500), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n206), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n523), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n504), .B2(new_n505), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n505), .A2(KEYINPUT30), .A3(new_n500), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT71), .A3(new_n206), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n522), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n520), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n534), .A2(new_n536), .A3(new_n521), .ZN(new_n537));
  INV_X1    g351(.A(new_n522), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT71), .B1(new_n532), .B2(new_n206), .ZN(new_n539));
  NOR4_X1   g353(.A1(new_n530), .A2(new_n531), .A3(new_n527), .A4(new_n509), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT73), .B1(new_n541), .B2(KEYINPUT31), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G472), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(KEYINPUT32), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n521), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n519), .B2(new_n515), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n536), .B1(new_n534), .B2(new_n521), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n541), .A2(KEYINPUT73), .A3(KEYINPUT31), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n544), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT76), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n519), .A2(KEYINPUT29), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n512), .A2(new_n493), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n505), .A2(new_n500), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n509), .A2(new_n510), .ZN(new_n560));
  AOI211_X1 g374(.A(KEYINPUT72), .B(new_n201), .C1(new_n226), .C2(new_n203), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n508), .A2(new_n511), .B1(new_n505), .B2(new_n500), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT74), .B(new_n558), .C1(new_n564), .C2(new_n493), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(KEYINPUT28), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n557), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n556), .B1(new_n568), .B2(new_n423), .ZN(new_n569));
  INV_X1    g383(.A(new_n563), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n493), .B1(new_n570), .B2(new_n512), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT76), .B(new_n356), .C1(new_n574), .C2(new_n557), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT29), .B1(new_n515), .B2(new_n519), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n562), .B1(new_n528), .B2(new_n533), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n519), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n543), .A2(KEYINPUT77), .A3(KEYINPUT32), .A4(new_n544), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n547), .A2(new_n555), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT24), .B(G110), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT80), .ZN(new_n584));
  XNOR2_X1  g398(.A(G119), .B(G128), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT23), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n194), .B2(G128), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n587), .B(new_n588), .C1(G119), .C2(new_n265), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n584), .A2(new_n585), .B1(G110), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n390), .A2(new_n391), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI22_X1  g406(.A1(new_n584), .A2(new_n585), .B1(G110), .B2(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(new_n380), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(G146), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n401), .A2(new_n406), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT22), .B(G137), .ZN(new_n598));
  INV_X1    g412(.A(G234), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n487), .A2(new_n599), .A3(G953), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n598), .B(new_n600), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n592), .B(new_n601), .C1(new_n595), .C2(new_n596), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT25), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n603), .A2(new_n356), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n349), .B1(new_n423), .B2(new_n599), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT79), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n603), .A2(new_n356), .A3(new_n604), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n605), .B2(KEYINPUT25), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n603), .A2(new_n604), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n609), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n492), .A2(new_n582), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(new_n617), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n491), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n551), .A2(new_n552), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n554), .B1(new_n622), .B2(new_n535), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n553), .B2(new_n423), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT101), .ZN(new_n627));
  INV_X1    g441(.A(new_n301), .ZN(new_n628));
  INV_X1    g442(.A(new_n371), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(new_n352), .B2(new_n336), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n355), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n633), .A2(KEYINPUT33), .A3(new_n354), .A4(new_n351), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n423), .A2(new_n357), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n355), .A2(new_n356), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n357), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n418), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n628), .A2(new_n629), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n627), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AOI21_X1  g459(.A(new_n418), .B1(new_n363), .B2(new_n365), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(new_n305), .A3(new_n187), .A4(new_n629), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n627), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND2_X1  g465(.A1(new_n543), .A2(new_n356), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n623), .B1(new_n652), .B2(G472), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n597), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n597), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n656), .A2(new_n615), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n610), .B2(new_n612), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n489), .B(new_n659), .C1(new_n477), .C2(new_n485), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n302), .A2(new_n307), .A3(new_n660), .A4(new_n419), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT37), .B(G110), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  INV_X1    g478(.A(new_n660), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n301), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n582), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n369), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n670));
  INV_X1    g484(.A(new_n368), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n646), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n305), .B(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n418), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n363), .B2(new_n365), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n187), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n673), .B(KEYINPUT39), .Z(new_n684));
  NAND3_X1  g498(.A1(new_n486), .A2(new_n490), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n519), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n577), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n564), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n279), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n547), .A2(new_n693), .A3(new_n555), .A4(new_n581), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n688), .A2(new_n659), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND2_X1  g510(.A1(new_n640), .A2(new_n674), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n667), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT105), .B(G146), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G48));
  AND2_X1   g515(.A1(new_n582), .A2(new_n617), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n471), .A2(new_n475), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(new_n423), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n476), .A2(new_n421), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT106), .B1(new_n706), .B2(new_n488), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  INV_X1    g522(.A(new_n488), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n704), .A2(new_n708), .A3(new_n709), .A4(new_n705), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n641), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n702), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n647), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n702), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NOR4_X1   g532(.A1(new_n366), .A2(new_n371), .A3(new_n418), .A4(new_n659), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n628), .A2(new_n719), .A3(new_n710), .A4(new_n707), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n582), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND3_X1  g536(.A1(new_n682), .A2(new_n187), .A3(new_n305), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n711), .A2(new_n723), .A3(new_n371), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n567), .B(new_n689), .C1(new_n571), .C2(new_n572), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n725), .B(new_n726), .C1(new_n534), .C2(new_n521), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n549), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n541), .A2(KEYINPUT31), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n725), .B1(new_n729), .B2(new_n726), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n544), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT108), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(new_n544), .C1(new_n728), .C2(new_n730), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n732), .A2(new_n625), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n735), .A3(new_n617), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NOR2_X1   g551(.A1(new_n711), .A2(new_n301), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n698), .ZN(new_n739));
  AOI22_X1  g553(.A1(KEYINPUT108), .A2(new_n731), .B1(new_n652), .B2(G472), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  INV_X1    g555(.A(new_n659), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n734), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n732), .A2(new_n625), .A3(new_n742), .A4(new_n734), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n739), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(G125), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G27));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  INV_X1    g563(.A(new_n705), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n478), .B1(new_n483), .B2(new_n470), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n421), .B1(new_n751), .B2(new_n279), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n709), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n303), .A2(new_n304), .A3(new_n187), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n697), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n582), .A2(new_n749), .A3(new_n617), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n555), .A2(new_n580), .A3(new_n545), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n617), .A3(new_n755), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT111), .B(G131), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G33));
  NOR3_X1   g576(.A1(new_n675), .A2(new_n753), .A3(new_n754), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n582), .A2(new_n763), .A3(new_n617), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n681), .A2(new_n639), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  AND3_X1   g581(.A1(new_n654), .A2(new_n742), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n754), .B1(new_n768), .B2(KEYINPUT44), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n481), .B2(new_n484), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n751), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n422), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT46), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n750), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n774), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n488), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n778), .A2(KEYINPUT112), .A3(new_n684), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT112), .B1(new_n778), .B2(new_n684), .ZN(new_n780));
  OAI221_X1 g594(.A(new_n769), .B1(KEYINPUT44), .B2(new_n768), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  OR2_X1    g596(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n582), .A2(new_n617), .A3(new_n697), .A4(new_n754), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  INV_X1    g602(.A(new_n739), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n582), .B(new_n666), .C1(new_n676), .C2(new_n698), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n723), .A2(new_n673), .A3(new_n753), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n694), .A2(new_n795), .A3(new_n659), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n796), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n798), .B2(new_n746), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n756), .A2(new_n759), .A3(new_n764), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n361), .A2(new_n362), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n681), .A2(new_n802), .A3(new_n674), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n665), .A2(new_n754), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n582), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n582), .A2(new_n804), .A3(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n743), .A2(new_n745), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n755), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n801), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n582), .A2(new_n720), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n653), .A2(new_n621), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n639), .A2(new_n418), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n639), .A2(new_n418), .A3(KEYINPUT113), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n418), .A2(new_n802), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n302), .A3(new_n307), .A4(new_n629), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n814), .A2(new_n821), .B1(new_n654), .B2(new_n661), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n582), .B(new_n617), .C1(new_n712), .C2(new_n716), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n618), .A3(new_n736), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n812), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n800), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n821), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n302), .A2(new_n307), .A3(new_n419), .A4(new_n660), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(new_n626), .B1(new_n829), .B2(new_n653), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n618), .A3(new_n721), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n824), .A2(new_n736), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n807), .A2(new_n808), .B1(new_n810), .B2(new_n755), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n801), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n797), .A2(new_n799), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n827), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n800), .A2(new_n826), .A3(KEYINPUT53), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n835), .B2(new_n836), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n783), .B(new_n784), .C1(new_n490), .C2(new_n706), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n617), .A2(new_n735), .A3(new_n368), .A4(new_n767), .ZN(new_n846));
  INV_X1    g660(.A(new_n754), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n711), .A2(new_n754), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n850), .A2(new_n694), .A3(new_n620), .A4(new_n671), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n639), .A2(new_n418), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n845), .A2(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n767), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n850), .A2(new_n854), .A3(new_n671), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n810), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n680), .A2(new_n711), .A3(new_n187), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT50), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n757), .A2(new_n617), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT48), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n367), .B(G953), .C1(new_n851), .C2(new_n640), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n846), .A2(new_n738), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n844), .A2(new_n862), .A3(new_n863), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(G952), .A2(G953), .ZN(new_n871));
  INV_X1    g685(.A(new_n680), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n706), .B(KEYINPUT49), .Z(new_n873));
  NAND3_X1  g687(.A1(new_n617), .A2(new_n490), .A3(new_n187), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n766), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n870), .A2(new_n871), .B1(new_n694), .B2(new_n876), .ZN(G75));
  XNOR2_X1  g691(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n256), .A2(new_n277), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n299), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n356), .B1(new_n840), .B2(new_n841), .ZN(new_n881));
  AOI211_X1 g695(.A(KEYINPUT56), .B(new_n880), .C1(new_n881), .C2(new_n189), .ZN(new_n882));
  INV_X1    g696(.A(new_n880), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n840), .A2(new_n841), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n423), .A3(new_n189), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n878), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n356), .B(new_n190), .C1(new_n840), .C2(new_n841), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n880), .B1(new_n889), .B2(KEYINPUT56), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n885), .A2(new_n886), .A3(new_n883), .ZN(new_n891));
  INV_X1    g705(.A(new_n878), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n367), .A2(G953), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT117), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n888), .A2(new_n893), .A3(new_n895), .ZN(G51));
  INV_X1    g710(.A(new_n895), .ZN(new_n897));
  INV_X1    g711(.A(new_n703), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT118), .B1(new_n884), .B2(KEYINPUT54), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n844), .B2(KEYINPUT118), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n422), .B(KEYINPUT57), .Z(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n881), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(new_n773), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n897), .B1(new_n902), .B2(new_n904), .ZN(G54));
  NAND3_X1  g719(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  INV_X1    g720(.A(new_n412), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n906), .A2(KEYINPUT119), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n895), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT119), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G60));
  AND2_X1   g725(.A1(new_n632), .A2(new_n634), .ZN(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n839), .B2(new_n843), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n912), .B(new_n915), .C1(new_n917), .C2(new_n899), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n839), .B2(new_n843), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n912), .ZN(new_n921));
  INV_X1    g735(.A(new_n843), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n842), .B1(new_n840), .B2(new_n841), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n912), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n895), .A2(new_n918), .A3(new_n921), .A4(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(new_n656), .A2(new_n657), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n884), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(KEYINPUT121), .A3(new_n895), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n895), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n614), .B1(new_n884), .B2(new_n931), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n933), .B(KEYINPUT61), .C1(new_n935), .C2(new_n936), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(G66));
  INV_X1    g754(.A(G224), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n370), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n833), .B2(G953), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n251), .B(new_n255), .C1(G898), .C2(new_n275), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  XNOR2_X1  g759(.A(new_n532), .B(KEYINPUT122), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n402), .A2(new_n403), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n723), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n864), .C1(new_n779), .C2(new_n780), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n792), .A2(new_n794), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n781), .A2(new_n787), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n801), .B(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n275), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n275), .A2(G900), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT124), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n948), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n948), .B(KEYINPUT123), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n695), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n685), .A2(new_n754), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n702), .A2(new_n820), .A3(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n781), .A2(new_n787), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(new_n275), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n958), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n467), .B2(new_n668), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G72));
  NAND3_X1  g785(.A1(new_n952), .A2(new_n833), .A3(new_n953), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  AND3_X1   g789(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n689), .B(new_n577), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n975), .B1(new_n967), .B2(new_n825), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n690), .ZN(new_n980));
  INV_X1    g794(.A(new_n975), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n577), .A2(new_n519), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(KEYINPUT127), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n534), .B1(new_n983), .B2(KEYINPUT127), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n897), .B1(new_n884), .B2(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n978), .A2(new_n980), .A3(new_n987), .ZN(G57));
endmodule


