

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U552 ( .A(KEYINPUT65), .B(n560), .Z(n674) );
  INV_X1 U553 ( .A(n717), .ZN(n736) );
  OR2_X1 U554 ( .A1(n742), .A2(n741), .ZN(n527) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n546) );
  NOR2_X2 U556 ( .A1(n577), .A2(n534), .ZN(G160) );
  NAND2_X1 U557 ( .A1(n720), .A2(n721), .ZN(n722) );
  XNOR2_X1 U558 ( .A(n712), .B(KEYINPUT64), .ZN(n735) );
  NAND2_X1 U559 ( .A1(n531), .A2(n529), .ZN(n528) );
  NAND2_X1 U560 ( .A1(n518), .A2(n719), .ZN(n529) );
  NAND2_X1 U561 ( .A1(n533), .A2(n532), .ZN(n531) );
  NOR2_X1 U562 ( .A1(n776), .A2(n765), .ZN(n766) );
  INV_X1 U563 ( .A(KEYINPUT33), .ZN(n540) );
  INV_X1 U564 ( .A(n959), .ZN(n539) );
  NOR2_X1 U565 ( .A1(n536), .A2(n780), .ZN(n782) );
  NAND2_X1 U566 ( .A1(n521), .A2(n815), .ZN(n543) );
  INV_X1 U567 ( .A(n722), .ZN(n533) );
  INV_X1 U568 ( .A(KEYINPUT28), .ZN(n727) );
  NAND2_X1 U569 ( .A1(n528), .A2(n723), .ZN(n724) );
  INV_X1 U570 ( .A(n735), .ZN(n717) );
  XNOR2_X1 U571 ( .A(n523), .B(KEYINPUT104), .ZN(n754) );
  NAND2_X1 U572 ( .A1(n526), .A2(n524), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n527), .B(KEYINPUT31), .ZN(n526) );
  AND2_X1 U574 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U575 ( .A1(G164), .A2(G1384), .ZN(n710) );
  AND2_X1 U576 ( .A1(n537), .A2(n538), .ZN(n536) );
  INV_X1 U577 ( .A(G2105), .ZN(n545) );
  AND2_X2 U578 ( .A1(n545), .A2(G2104), .ZN(n567) );
  NAND2_X1 U579 ( .A1(n542), .A2(n832), .ZN(n541) );
  OR2_X1 U580 ( .A1(n783), .A2(n543), .ZN(n542) );
  XNOR2_X1 U581 ( .A(n535), .B(n573), .ZN(n534) );
  AND2_X1 U582 ( .A1(n718), .A2(n530), .ZN(n518) );
  OR2_X1 U583 ( .A1(n740), .A2(G301), .ZN(n519) );
  NAND2_X1 U584 ( .A1(n767), .A2(n766), .ZN(n520) );
  INV_X1 U585 ( .A(n958), .ZN(n532) );
  XOR2_X1 U586 ( .A(n709), .B(KEYINPUT93), .Z(n521) );
  XNOR2_X1 U587 ( .A(KEYINPUT103), .B(KEYINPUT29), .ZN(n522) );
  NAND2_X1 U588 ( .A1(n525), .A2(n519), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n731), .B(n522), .ZN(n525) );
  INV_X1 U590 ( .A(n955), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n711), .A2(G160), .ZN(n712) );
  NAND2_X1 U592 ( .A1(n571), .A2(n572), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n520), .A2(n540), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n769), .A2(n539), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n541), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X2 U596 ( .A(KEYINPUT17), .B(n546), .Z(n866) );
  AND2_X1 U597 ( .A1(n600), .A2(n599), .ZN(n544) );
  INV_X1 U598 ( .A(n945), .ZN(n762) );
  INV_X1 U599 ( .A(n946), .ZN(n765) );
  XNOR2_X1 U600 ( .A(n752), .B(KEYINPUT32), .ZN(n760) );
  INV_X1 U601 ( .A(KEYINPUT109), .ZN(n781) );
  AND2_X1 U602 ( .A1(n544), .A2(n605), .ZN(n606) );
  XOR2_X1 U603 ( .A(KEYINPUT1), .B(n558), .Z(n666) );
  NOR2_X1 U604 ( .A1(n552), .A2(n551), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G102), .A2(n567), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G138), .A2(n866), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n552) );
  AND2_X1 U608 ( .A1(G2104), .A2(G2105), .ZN(n862) );
  NAND2_X1 U609 ( .A1(G114), .A2(n862), .ZN(n550) );
  NOR2_X1 U610 ( .A1(G2104), .A2(n545), .ZN(n863) );
  NAND2_X1 U611 ( .A1(G126), .A2(n863), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U613 ( .A1(G651), .A2(G543), .ZN(n667) );
  NAND2_X1 U614 ( .A1(n667), .A2(G89), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  INV_X1 U617 ( .A(G651), .ZN(n557) );
  NOR2_X1 U618 ( .A1(n650), .A2(n557), .ZN(n670) );
  NAND2_X1 U619 ( .A1(G76), .A2(n670), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT5), .ZN(n565) );
  NOR2_X1 U622 ( .A1(G543), .A2(n557), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n666), .A2(G63), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT76), .ZN(n562) );
  NOR2_X1 U625 ( .A1(G651), .A2(n650), .ZN(n560) );
  NAND2_X1 U626 ( .A1(G51), .A2(n674), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U632 ( .A(KEYINPUT67), .ZN(n573) );
  INV_X1 U633 ( .A(KEYINPUT23), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G101), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT66), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G125), .A2(n863), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G137), .A2(n866), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G113), .A2(n862), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT68), .B(n576), .ZN(n577) );
  AND2_X1 U642 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U643 ( .A(G132), .ZN(G219) );
  INV_X1 U644 ( .A(G82), .ZN(G220) );
  NAND2_X1 U645 ( .A1(G64), .A2(n666), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G52), .A2(n674), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G90), .A2(n667), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G77), .A2(n670), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT9), .B(n582), .Z(n583) );
  NOR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(G171) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n833) );
  NAND2_X1 U656 ( .A1(n833), .A2(G567), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n586), .B(KEYINPUT71), .ZN(n587) );
  XNOR2_X1 U658 ( .A(KEYINPUT11), .B(n587), .ZN(G234) );
  XOR2_X1 U659 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n589) );
  NAND2_X1 U660 ( .A1(G56), .A2(n666), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n589), .B(n588), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n667), .A2(G81), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G68), .A2(n670), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT13), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G43), .A2(n674), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U670 ( .A(KEYINPUT73), .B(n598), .ZN(n955) );
  INV_X1 U671 ( .A(G860), .ZN(n619) );
  OR2_X1 U672 ( .A1(n955), .A2(n619), .ZN(G153) );
  INV_X1 U673 ( .A(G171), .ZN(G301) );
  NAND2_X1 U674 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G79), .A2(n670), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G54), .A2(n674), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n667), .A2(G92), .ZN(n601) );
  XNOR2_X1 U678 ( .A(n601), .B(KEYINPUT74), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G66), .A2(n666), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT75), .ZN(n605) );
  XNOR2_X1 U682 ( .A(KEYINPUT15), .B(n606), .ZN(n958) );
  INV_X1 U683 ( .A(G868), .ZN(n687) );
  NAND2_X1 U684 ( .A1(n958), .A2(n687), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G284) );
  NAND2_X1 U686 ( .A1(G65), .A2(n666), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G91), .A2(n667), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G78), .A2(n670), .ZN(n611) );
  XNOR2_X1 U690 ( .A(KEYINPUT69), .B(n611), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n674), .A2(G53), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G299) );
  NOR2_X1 U694 ( .A1(G286), .A2(n687), .ZN(n616) );
  XOR2_X1 U695 ( .A(KEYINPUT77), .B(n616), .Z(n618) );
  NOR2_X1 U696 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G297) );
  NAND2_X1 U698 ( .A1(n619), .A2(G559), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n620), .A2(n532), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n621), .B(KEYINPUT16), .ZN(n622) );
  XNOR2_X1 U701 ( .A(KEYINPUT78), .B(n622), .ZN(G148) );
  NOR2_X1 U702 ( .A1(G559), .A2(n687), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n532), .A2(n623), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n624), .B(KEYINPUT79), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n955), .A2(G868), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT80), .B(n627), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G99), .A2(n567), .ZN(n628) );
  XOR2_X1 U709 ( .A(KEYINPUT82), .B(n628), .Z(n634) );
  NAND2_X1 U710 ( .A1(n863), .A2(G123), .ZN(n629) );
  XNOR2_X1 U711 ( .A(n629), .B(KEYINPUT18), .ZN(n631) );
  NAND2_X1 U712 ( .A1(G135), .A2(n866), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U714 ( .A(KEYINPUT81), .B(n632), .Z(n633) );
  NOR2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n862), .A2(G111), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n1007) );
  XNOR2_X1 U718 ( .A(G2096), .B(n1007), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n637), .A2(G2100), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(KEYINPUT83), .ZN(G156) );
  NAND2_X1 U721 ( .A1(G559), .A2(n532), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n639), .B(n955), .ZN(n684) );
  NOR2_X1 U723 ( .A1(n684), .A2(G860), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G67), .A2(n666), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G93), .A2(n667), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G80), .A2(n670), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G55), .A2(n674), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n644) );
  OR2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n688) );
  XOR2_X1 U731 ( .A(n646), .B(n688), .Z(G145) );
  NAND2_X1 U732 ( .A1(G49), .A2(n674), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U735 ( .A1(n666), .A2(n649), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G288) );
  AND2_X1 U738 ( .A1(n666), .A2(G60), .ZN(n656) );
  NAND2_X1 U739 ( .A1(G85), .A2(n667), .ZN(n654) );
  NAND2_X1 U740 ( .A1(G72), .A2(n670), .ZN(n653) );
  NAND2_X1 U741 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U742 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U743 ( .A1(n674), .A2(G47), .ZN(n657) );
  NAND2_X1 U744 ( .A1(n658), .A2(n657), .ZN(G290) );
  NAND2_X1 U745 ( .A1(G62), .A2(n666), .ZN(n660) );
  NAND2_X1 U746 ( .A1(G88), .A2(n667), .ZN(n659) );
  NAND2_X1 U747 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n670), .A2(G75), .ZN(n661) );
  XOR2_X1 U749 ( .A(KEYINPUT84), .B(n661), .Z(n662) );
  NOR2_X1 U750 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n674), .A2(G50), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n665), .A2(n664), .ZN(G303) );
  NAND2_X1 U753 ( .A1(G61), .A2(n666), .ZN(n669) );
  NAND2_X1 U754 ( .A1(G86), .A2(n667), .ZN(n668) );
  NAND2_X1 U755 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U756 ( .A1(n670), .A2(G73), .ZN(n671) );
  XOR2_X1 U757 ( .A(KEYINPUT2), .B(n671), .Z(n672) );
  NOR2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n674), .A2(G48), .ZN(n675) );
  NAND2_X1 U760 ( .A1(n676), .A2(n675), .ZN(G305) );
  XNOR2_X1 U761 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n678) );
  XNOR2_X1 U762 ( .A(G288), .B(KEYINPUT19), .ZN(n677) );
  XNOR2_X1 U763 ( .A(n678), .B(n677), .ZN(n679) );
  XOR2_X1 U764 ( .A(n688), .B(n679), .Z(n681) );
  INV_X1 U765 ( .A(G299), .ZN(n948) );
  XNOR2_X1 U766 ( .A(G290), .B(n948), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n682), .B(G303), .ZN(n683) );
  XNOR2_X1 U769 ( .A(n683), .B(G305), .ZN(n889) );
  XNOR2_X1 U770 ( .A(n889), .B(n684), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n685), .A2(G868), .ZN(n686) );
  XOR2_X1 U772 ( .A(KEYINPUT87), .B(n686), .Z(n690) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n690), .A2(n689), .ZN(G295) );
  NAND2_X1 U775 ( .A1(G2078), .A2(G2084), .ZN(n691) );
  XOR2_X1 U776 ( .A(KEYINPUT20), .B(n691), .Z(n692) );
  NAND2_X1 U777 ( .A1(G2090), .A2(n692), .ZN(n695) );
  XOR2_X1 U778 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n693) );
  XNOR2_X1 U779 ( .A(KEYINPUT21), .B(n693), .ZN(n694) );
  XNOR2_X1 U780 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U781 ( .A1(n696), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U782 ( .A(n697), .B(KEYINPUT90), .ZN(G158) );
  XOR2_X1 U783 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XOR2_X1 U784 ( .A(KEYINPUT91), .B(G44), .Z(n698) );
  XNOR2_X1 U785 ( .A(KEYINPUT3), .B(n698), .ZN(G218) );
  NAND2_X1 U786 ( .A1(G483), .A2(G661), .ZN(n706) );
  NAND2_X1 U787 ( .A1(G108), .A2(G120), .ZN(n699) );
  NOR2_X1 U788 ( .A1(G237), .A2(n699), .ZN(n700) );
  NAND2_X1 U789 ( .A1(G69), .A2(n700), .ZN(n837) );
  NAND2_X1 U790 ( .A1(n837), .A2(G567), .ZN(n705) );
  NOR2_X1 U791 ( .A1(G220), .A2(G219), .ZN(n701) );
  XOR2_X1 U792 ( .A(KEYINPUT22), .B(n701), .Z(n702) );
  NOR2_X1 U793 ( .A1(G218), .A2(n702), .ZN(n703) );
  NAND2_X1 U794 ( .A1(G96), .A2(n703), .ZN(n838) );
  NAND2_X1 U795 ( .A1(n838), .A2(G2106), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n918) );
  NOR2_X1 U797 ( .A1(n706), .A2(n918), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n707), .B(KEYINPUT92), .ZN(n836) );
  NAND2_X1 U799 ( .A1(G36), .A2(n836), .ZN(G176) );
  INV_X1 U800 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U801 ( .A(G1986), .B(G290), .ZN(n944) );
  NAND2_X1 U802 ( .A1(G160), .A2(G40), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n710), .A2(n708), .ZN(n829) );
  NAND2_X1 U804 ( .A1(n944), .A2(n829), .ZN(n709) );
  AND2_X1 U805 ( .A1(n710), .A2(G40), .ZN(n711) );
  NAND2_X1 U806 ( .A1(G2072), .A2(n717), .ZN(n713) );
  XNOR2_X1 U807 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  INV_X1 U808 ( .A(G1956), .ZN(n919) );
  NOR2_X1 U809 ( .A1(n717), .A2(n919), .ZN(n714) );
  NOR2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n726) );
  NAND2_X1 U811 ( .A1(n948), .A2(n726), .ZN(n725) );
  NAND2_X1 U812 ( .A1(n717), .A2(G1996), .ZN(n716) );
  XNOR2_X1 U813 ( .A(n716), .B(KEYINPUT26), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n736), .A2(G1341), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n736), .A2(G1348), .ZN(n721) );
  NAND2_X1 U816 ( .A1(G2067), .A2(n717), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n958), .A2(n722), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n948), .A2(n726), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U822 ( .A(KEYINPUT25), .B(G2078), .Z(n976) );
  NOR2_X1 U823 ( .A1(n736), .A2(n976), .ZN(n732) );
  XNOR2_X1 U824 ( .A(n732), .B(KEYINPUT102), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n717), .A2(G1961), .ZN(n733) );
  NOR2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n735), .A2(G8), .ZN(n776) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n776), .ZN(n756) );
  NOR2_X1 U829 ( .A1(n736), .A2(G2084), .ZN(n753) );
  NOR2_X1 U830 ( .A1(n756), .A2(n753), .ZN(n737) );
  NAND2_X1 U831 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U832 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U833 ( .A1(G168), .A2(n739), .ZN(n742) );
  AND2_X1 U834 ( .A1(G301), .A2(n740), .ZN(n741) );
  NAND2_X1 U835 ( .A1(n754), .A2(G286), .ZN(n750) );
  NOR2_X1 U836 ( .A1(n736), .A2(G2090), .ZN(n743) );
  XOR2_X1 U837 ( .A(KEYINPUT105), .B(n743), .Z(n745) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n776), .ZN(n744) );
  NOR2_X1 U839 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U840 ( .A(KEYINPUT106), .B(n746), .Z(n747) );
  NOR2_X1 U841 ( .A1(G166), .A2(n747), .ZN(n748) );
  XNOR2_X1 U842 ( .A(n748), .B(KEYINPUT107), .ZN(n749) );
  NAND2_X1 U843 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n751), .A2(G8), .ZN(n752) );
  NAND2_X1 U845 ( .A1(G8), .A2(n753), .ZN(n758) );
  INV_X1 U846 ( .A(n754), .ZN(n755) );
  NOR2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n770) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n761) );
  XOR2_X1 U851 ( .A(n761), .B(KEYINPUT108), .Z(n763) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n945) );
  NAND2_X1 U853 ( .A1(n770), .A2(n764), .ZN(n767) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n946) );
  NAND2_X1 U855 ( .A1(n945), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n768), .A2(n776), .ZN(n769) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n959) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n770), .A2(n772), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n776), .A2(n773), .ZN(n779) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT24), .ZN(n775) );
  XNOR2_X1 U864 ( .A(n775), .B(KEYINPUT101), .ZN(n777) );
  OR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n782), .B(n781), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G95), .A2(n567), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G131), .A2(n866), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U871 ( .A1(G119), .A2(n863), .ZN(n786) );
  XNOR2_X1 U872 ( .A(KEYINPUT97), .B(n786), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n862), .A2(G107), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n850) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n850), .ZN(n791) );
  XNOR2_X1 U877 ( .A(n791), .B(KEYINPUT98), .ZN(n801) );
  NAND2_X1 U878 ( .A1(G117), .A2(n862), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G129), .A2(n863), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n567), .A2(G105), .ZN(n794) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n794), .Z(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U884 ( .A(KEYINPUT99), .B(n797), .Z(n799) );
  NAND2_X1 U885 ( .A1(n866), .A2(G141), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n846) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n846), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U889 ( .A(KEYINPUT100), .B(n802), .ZN(n1006) );
  NAND2_X1 U890 ( .A1(n829), .A2(n1006), .ZN(n817) );
  XNOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  XNOR2_X1 U892 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G104), .A2(n567), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G140), .A2(n866), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U896 ( .A(n806), .B(n805), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G128), .A2(n863), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n862), .A2(G116), .ZN(n807) );
  XOR2_X1 U899 ( .A(KEYINPUT95), .B(n807), .Z(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n810), .B(KEYINPUT96), .ZN(n811) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n811), .Z(n812) );
  NOR2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n814), .ZN(n874) );
  NOR2_X1 U905 ( .A1(n827), .A2(n874), .ZN(n1001) );
  NAND2_X1 U906 ( .A1(n1001), .A2(n829), .ZN(n816) );
  AND2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n815) );
  INV_X1 U908 ( .A(n816), .ZN(n826) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n846), .ZN(n1003) );
  INV_X1 U910 ( .A(n817), .ZN(n820) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n850), .ZN(n1010) );
  NOR2_X1 U913 ( .A1(n818), .A2(n1010), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n1003), .A2(n821), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT39), .ZN(n823) );
  XNOR2_X1 U917 ( .A(KEYINPUT110), .B(n823), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(n829), .ZN(n825) );
  OR2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n874), .A2(n827), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n828), .B(KEYINPUT111), .ZN(n1015) );
  NAND2_X1 U922 ( .A1(n1015), .A2(n829), .ZN(n830) );
  AND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U926 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  NAND2_X1 U936 ( .A1(G124), .A2(n863), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(KEYINPUT44), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n567), .A2(G100), .ZN(n840) );
  NAND2_X1 U939 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U940 ( .A1(G136), .A2(n866), .ZN(n843) );
  NAND2_X1 U941 ( .A1(G112), .A2(n862), .ZN(n842) );
  NAND2_X1 U942 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U943 ( .A1(n845), .A2(n844), .ZN(G162) );
  XNOR2_X1 U944 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n846), .B(KEYINPUT115), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G160), .B(G162), .Z(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(n861) );
  NAND2_X1 U950 ( .A1(G103), .A2(n567), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G139), .A2(n866), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U953 ( .A1(G115), .A2(n862), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G127), .A2(n863), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n996) );
  XNOR2_X1 U958 ( .A(G164), .B(n996), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n876) );
  NAND2_X1 U960 ( .A1(G118), .A2(n862), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G130), .A2(n863), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U963 ( .A1(G106), .A2(n567), .ZN(n868) );
  NAND2_X1 U964 ( .A1(G142), .A2(n866), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U966 ( .A(n869), .B(KEYINPUT45), .Z(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(n1007), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U970 ( .A(n876), .B(n875), .ZN(n877) );
  NOR2_X1 U971 ( .A1(G37), .A2(n877), .ZN(G395) );
  XNOR2_X1 U972 ( .A(G2454), .B(G2451), .ZN(n886) );
  XNOR2_X1 U973 ( .A(G2430), .B(G2446), .ZN(n884) );
  XOR2_X1 U974 ( .A(G2435), .B(G2427), .Z(n879) );
  XNOR2_X1 U975 ( .A(KEYINPUT112), .B(G2438), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U977 ( .A(n880), .B(G2443), .Z(n882) );
  XNOR2_X1 U978 ( .A(G1341), .B(G1348), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n887) );
  NAND2_X1 U982 ( .A1(n887), .A2(G14), .ZN(n888) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(n888), .ZN(G401) );
  XNOR2_X1 U984 ( .A(G286), .B(n889), .ZN(n891) );
  XNOR2_X1 U985 ( .A(n958), .B(G171), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n892), .B(n955), .ZN(n893) );
  NOR2_X1 U988 ( .A1(G37), .A2(n893), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2100), .B(G2096), .Z(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT42), .B(G2678), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U992 ( .A(KEYINPUT43), .B(G2090), .Z(n897) );
  XNOR2_X1 U993 ( .A(G2067), .B(G2072), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U996 ( .A(G2078), .B(G2084), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(G227) );
  XNOR2_X1 U998 ( .A(G1996), .B(KEYINPUT114), .ZN(n911) );
  XOR2_X1 U999 ( .A(G1976), .B(G1971), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G1991), .B(G1986), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1002 ( .A(G1981), .B(G1961), .Z(n905) );
  XNOR2_X1 U1003 ( .A(G1966), .B(G1956), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1006 ( .A(G2474), .B(KEYINPUT41), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(G229) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n918), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(G397), .A2(n913), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(n916), .ZN(n917) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(n917), .Z(G225) );
  XNOR2_X1 U1016 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n918), .ZN(G319) );
  XNOR2_X1 U1018 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1024) );
  XOR2_X1 U1019 ( .A(G1966), .B(G21), .Z(n930) );
  XNOR2_X1 U1020 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(G20), .B(n919), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(G1341), .B(G19), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(G1981), .B(G6), .ZN(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n926) );
  XOR2_X1 U1026 ( .A(KEYINPUT59), .B(G1348), .Z(n924) );
  XNOR2_X1 U1027 ( .A(G4), .B(n924), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(n928), .B(n927), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT125), .B(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G1961), .B(G5), .Z(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G22), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(G23), .B(G1976), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1037 ( .A(G1986), .B(G24), .Z(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(n938), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n941), .Z(n942) );
  NOR2_X1 U1042 ( .A1(G16), .A2(n942), .ZN(n994) );
  XNOR2_X1 U1043 ( .A(KEYINPUT56), .B(G16), .ZN(n968) );
  XNOR2_X1 U1044 ( .A(G1961), .B(G171), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(n943), .B(KEYINPUT122), .ZN(n954) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G166), .B(G1971), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n948), .B(G1956), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(n958), .B(G1348), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(n961), .B(KEYINPUT57), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(KEYINPUT121), .B(n962), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT123), .ZN(n991) );
  XNOR2_X1 U1064 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n988) );
  XNOR2_X1 U1065 ( .A(G2084), .B(G34), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n970), .B(KEYINPUT54), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G35), .B(G2090), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n986) );
  XOR2_X1 U1069 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n984) );
  XOR2_X1 U1070 ( .A(G1991), .B(G25), .Z(n973) );
  NAND2_X1 U1071 ( .A1(n973), .A2(G28), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G32), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(G33), .B(G2072), .ZN(n974) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(G2067), .B(G26), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(G27), .B(n976), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1080 ( .A(n984), .B(n983), .Z(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n988), .B(n987), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n989), .A2(G29), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(G11), .A2(n992), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT126), .ZN(n1022) );
  XOR2_X1 U1088 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1091 ( .A(KEYINPUT50), .B(n999), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1017) );
  XOR2_X1 U1093 ( .A(G2090), .B(G162), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(KEYINPUT51), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT118), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1018), .ZN(n1019) );
  OR2_X1 U1105 ( .A1(KEYINPUT55), .A2(n1019), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(G29), .A2(n1020), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1024), .B(n1023), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

