//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n203), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT64), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n201), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n203), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n247), .B(new_n252), .ZN(G351));
  AND2_X1   g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT5), .A2(G41), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT5), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(G270), .B(new_n256), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n254), .B2(new_n255), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT5), .B(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n256), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n273), .A3(G257), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G303), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n274), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n271), .A2(new_n273), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n231), .A3(new_n275), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n269), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n268), .A2(new_n285), .A3(G179), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT83), .A2(G116), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT83), .A2(G116), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G283), .ZN(new_n291));
  INV_X1    g0091(.A(G97), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n291), .B(new_n210), .C1(G33), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n219), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n290), .A2(KEYINPUT20), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n295), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n287), .A2(new_n288), .A3(new_n210), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n209), .A2(G33), .ZN(new_n303));
  AND4_X1   g0103(.A1(new_n219), .A2(new_n302), .A3(new_n294), .A4(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n302), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n304), .A2(G116), .B1(new_n305), .B2(new_n289), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n301), .A2(KEYINPUT86), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT86), .B1(new_n301), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n286), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n286), .B(KEYINPUT87), .C1(new_n307), .C2(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n307), .A2(new_n308), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n268), .A2(new_n285), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n314), .B(new_n316), .C1(new_n317), .C2(new_n315), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT21), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n268), .A2(new_n285), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G169), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(KEYINPUT21), .C1(new_n308), .C2(new_n307), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n313), .A2(new_n318), .A3(new_n322), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT88), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n322), .A2(new_n325), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n329), .A2(KEYINPUT88), .A3(new_n313), .A4(new_n318), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G294), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT66), .B(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n280), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n332), .B1(new_n334), .B2(new_n225), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n274), .A2(new_n275), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n269), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n256), .B1(new_n259), .B2(new_n262), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G264), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n267), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n267), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n323), .ZN(new_n345));
  INV_X1    g0145(.A(new_n295), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT24), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n280), .A2(new_n210), .A3(G87), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT22), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT22), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n280), .A2(new_n350), .A3(new_n210), .A4(G87), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n289), .A2(new_n270), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT23), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n210), .B2(G107), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n353), .A2(new_n210), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n347), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n347), .A3(new_n357), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n346), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT25), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n302), .B2(G107), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n302), .A2(new_n362), .A3(G107), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n363), .A2(new_n365), .B1(new_n304), .B2(G107), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n343), .B(new_n345), .C1(new_n361), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n352), .A2(new_n347), .A3(new_n357), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n295), .B1(new_n370), .B2(new_n358), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n344), .A2(G200), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n337), .A2(G190), .A3(new_n267), .A4(new_n340), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n366), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT85), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n280), .A2(new_n333), .A3(G244), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n280), .A2(new_n333), .A3(KEYINPUT4), .A4(G244), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n381), .A2(new_n291), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n269), .ZN(new_n385));
  INV_X1    g0185(.A(G257), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n267), .B1(new_n338), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n378), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  AOI211_X1 g0189(.A(KEYINPUT80), .B(new_n387), .C1(new_n384), .C2(new_n269), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n323), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(new_n388), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(KEYINPUT67), .A2(G179), .ZN(new_n394));
  NOR2_X1   g0194(.A1(KEYINPUT67), .A2(G179), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n302), .A2(G97), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n304), .B2(G97), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT79), .ZN(new_n402));
  NAND2_X1  g0202(.A1(KEYINPUT6), .A2(G107), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT77), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(KEYINPUT6), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G97), .A2(G107), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n207), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n406), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n408), .A2(new_n206), .B1(new_n404), .B2(KEYINPUT6), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT78), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n210), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(G20), .A2(G33), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(new_n228), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n402), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n280), .B2(G20), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT73), .B(new_n419), .C1(new_n280), .C2(G20), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(G107), .A3(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n407), .A2(new_n412), .A3(new_n409), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n412), .B1(new_n407), .B2(new_n409), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n417), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(KEYINPUT79), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n418), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n401), .B1(new_n431), .B2(new_n295), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n398), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n425), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT79), .B1(new_n428), .B2(new_n429), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n295), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n383), .A2(new_n291), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n380), .B2(new_n379), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n256), .B1(new_n438), .B2(new_n382), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT80), .B1(new_n439), .B2(new_n387), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n385), .A2(new_n378), .A3(new_n388), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(G190), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n392), .A2(G200), .ZN(new_n443));
  AND4_X1   g0243(.A1(new_n436), .A2(new_n400), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT81), .B1(new_n433), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n441), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n323), .B1(new_n396), .B2(new_n393), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(new_n400), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT81), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n436), .A2(new_n400), .A3(new_n442), .A4(new_n443), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT15), .B(G87), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n302), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n280), .A2(new_n210), .A3(G68), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT19), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n210), .A2(G33), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(new_n292), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G97), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n210), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n206), .A2(new_n224), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT84), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n456), .B(new_n459), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n455), .B1(new_n465), .B2(new_n295), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n346), .A2(new_n302), .A3(new_n303), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n466), .B1(new_n453), .B2(new_n467), .ZN(new_n468));
  AND4_X1   g0268(.A1(new_n271), .A2(new_n273), .A3(new_n276), .A4(new_n278), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n353), .B1(G238), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n229), .A2(new_n275), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n280), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT82), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n280), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n256), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n269), .A2(new_n261), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G250), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n265), .A2(new_n261), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n323), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n475), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n474), .B1(new_n280), .B2(new_n471), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n334), .A2(new_n223), .B1(new_n270), .B2(new_n289), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n269), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n481), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(new_n396), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n468), .A2(new_n482), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(G200), .B1(new_n477), .B2(new_n481), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n488), .A3(G190), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n467), .A2(new_n224), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n455), .B(new_n493), .C1(new_n465), .C2(new_n295), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AND4_X1   g0297(.A1(new_n377), .A2(new_n445), .A3(new_n452), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n451), .B1(new_n432), .B2(new_n398), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(KEYINPUT81), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n377), .B1(new_n500), .B2(new_n452), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n331), .B(new_n376), .C1(new_n498), .C2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT65), .ZN(new_n503));
  INV_X1    g0303(.A(G41), .ZN(new_n504));
  AOI21_X1  g0304(.A(G1), .B1(new_n504), .B2(new_n260), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n503), .B1(new_n265), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n265), .A2(new_n503), .A3(new_n505), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n269), .A2(new_n505), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n507), .A2(new_n508), .B1(G238), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G226), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n460), .B1(new_n334), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G232), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n283), .A2(new_n513), .A3(new_n275), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n269), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT13), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT13), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n510), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  OR3_X1    g0321(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n305), .A2(new_n295), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n209), .A2(G20), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G68), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n458), .A2(new_n228), .B1(new_n210), .B2(G68), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT70), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(new_n201), .B2(new_n416), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n295), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT11), .ZN(new_n534));
  OAI221_X1 g0334(.A(new_n524), .B1(new_n526), .B2(new_n528), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n517), .A2(G190), .A3(new_n519), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n521), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT71), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n521), .A2(new_n537), .A3(KEYINPUT71), .A4(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n283), .A2(new_n275), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(G223), .B1(G77), .B2(new_n283), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n469), .A2(G222), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n256), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n265), .A2(new_n503), .A3(new_n505), .ZN(new_n548));
  INV_X1    g0348(.A(new_n505), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n256), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n548), .A2(new_n506), .B1(new_n511), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n396), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n552), .A2(G169), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT8), .B(G58), .ZN(new_n557));
  INV_X1    g0357(.A(G150), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n557), .A2(new_n458), .B1(new_n558), .B2(new_n416), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G20), .B2(new_n204), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n346), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n201), .B1(new_n209), .B2(G20), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n525), .A2(new_n562), .B1(new_n201), .B2(new_n305), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n555), .A2(new_n556), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT9), .B1(new_n561), .B2(new_n564), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n563), .C1(new_n560), .C2(new_n346), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n567), .A2(new_n569), .B1(new_n552), .B2(G190), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT69), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n553), .A2(new_n571), .A3(G200), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT69), .B1(new_n552), .B2(new_n317), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT10), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT10), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n570), .A2(new_n572), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n566), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n537), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT14), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n520), .A2(new_n580), .A3(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n342), .B2(new_n520), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n580), .B1(new_n520), .B2(G169), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n544), .A2(G238), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n230), .B2(new_n280), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n283), .A2(new_n279), .A3(new_n513), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n269), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n507), .A2(new_n508), .B1(G244), .B2(new_n509), .ZN(new_n589));
  AOI21_X1  g0389(.A(G169), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n557), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(new_n415), .B1(G20), .B2(G77), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n458), .B2(new_n453), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n593), .A2(new_n295), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n525), .A2(G77), .A3(new_n527), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G77), .B2(new_n302), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n588), .A2(new_n589), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(KEYINPUT68), .B1(new_n396), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT68), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n590), .B2(new_n597), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n588), .A2(new_n589), .ZN(new_n603));
  AOI211_X1 g0403(.A(new_n594), .B(new_n596), .C1(new_n603), .C2(G200), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(G190), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n600), .A2(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n543), .A2(new_n578), .A3(new_n584), .A4(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(G1698), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT74), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT74), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n280), .A2(new_n610), .A3(G226), .A4(G1698), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G223), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n334), .A2(new_n613), .B1(new_n270), .B2(new_n224), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n269), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n548), .A2(new_n506), .B1(new_n513), .B2(new_n550), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n323), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n270), .A2(new_n224), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n469), .B2(G223), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(new_n611), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n256), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n622), .A2(new_n616), .A3(new_n396), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT75), .B1(new_n618), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(new_n617), .A3(new_n554), .ZN(new_n625));
  OAI21_X1  g0425(.A(G169), .B1(new_n622), .B2(new_n616), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT75), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n591), .A2(new_n527), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n526), .A2(new_n630), .B1(new_n302), .B2(new_n591), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n423), .A2(G68), .A3(new_n424), .ZN(new_n632));
  XNOR2_X1  g0432(.A(G58), .B(G68), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(G20), .B1(G159), .B2(new_n415), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT16), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n346), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT72), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n420), .A2(new_n421), .A3(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n283), .A2(KEYINPUT72), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G68), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT16), .A3(new_n634), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT18), .B1(new_n629), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n317), .B1(new_n615), .B2(new_n617), .ZN(new_n645));
  INV_X1    g0445(.A(G190), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n622), .A2(new_n616), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT17), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n635), .A2(new_n636), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n295), .A3(new_n642), .ZN(new_n653));
  INV_X1    g0453(.A(new_n631), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT18), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n624), .A4(new_n628), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n643), .A2(KEYINPUT17), .A3(new_n648), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n644), .A2(new_n651), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT76), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT76), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n607), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n502), .A2(new_n664), .ZN(G372));
  NAND2_X1  g0465(.A1(new_n575), .A2(new_n577), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n651), .A2(new_n658), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n600), .A2(new_n602), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n543), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n669), .B2(new_n584), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n644), .A2(new_n657), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n566), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n664), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n313), .A2(new_n368), .A3(new_n322), .A4(new_n325), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n375), .A2(new_n496), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n449), .A3(new_n451), .A4(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT26), .B1(new_n433), .B2(new_n497), .ZN(new_n680));
  AND4_X1   g0480(.A1(KEYINPUT26), .A2(new_n497), .A3(new_n447), .A4(new_n448), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n679), .B(new_n490), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(G369));
  NAND2_X1  g0484(.A1(new_n329), .A2(new_n313), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n688), .A3(G213), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n314), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n693), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n331), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT89), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(G330), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT89), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n692), .B1(new_n371), .B2(new_n366), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n368), .B1(new_n375), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n368), .B2(new_n691), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n685), .A2(new_n692), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n705), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n369), .B2(new_n692), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n213), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n462), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n217), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n331), .A2(new_n376), .A3(new_n692), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n498), .B2(new_n501), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n477), .A2(new_n481), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n721), .A2(new_n286), .A3(new_n341), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n389), .A2(new_n390), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT30), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n721), .A2(new_n554), .A3(new_n315), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n344), .A3(new_n392), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n691), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n700), .B1(new_n720), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n682), .B2(new_n692), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n682), .A2(new_n735), .A3(new_n692), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n718), .B1(new_n740), .B2(G1), .ZN(G364));
  AND2_X1   g0541(.A1(new_n210), .A2(G13), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G1), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n713), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT90), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT90), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n213), .A2(G355), .A3(new_n280), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n712), .A2(new_n280), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G45), .B2(new_n217), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n252), .A2(new_n260), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(G116), .B2(new_n213), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n219), .B1(G20), .B2(new_n323), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n748), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n317), .A2(G179), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n210), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G283), .A2(new_n764), .B1(new_n767), .B2(G329), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n210), .A2(new_n646), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n761), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n768), .B(new_n283), .C1(new_n281), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n554), .A2(new_n317), .A3(new_n769), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n210), .A2(new_n317), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n554), .A2(new_n646), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G322), .A2(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n554), .A2(G190), .A3(new_n774), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n554), .A2(new_n317), .A3(new_n762), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G326), .A2(new_n780), .B1(new_n782), .B2(G311), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n765), .A2(G190), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n771), .B(new_n784), .C1(G294), .C2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G50), .A2(new_n780), .B1(new_n773), .B2(G58), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n228), .B2(new_n781), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  INV_X1    g0590(.A(new_n770), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n283), .B1(new_n791), .B2(G87), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n792), .A2(KEYINPUT92), .B1(new_n203), .B2(new_n775), .ZN(new_n793));
  INV_X1    g0593(.A(new_n786), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n292), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n764), .A2(G107), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  OR3_X1    g0598(.A1(new_n766), .A2(KEYINPUT32), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(KEYINPUT32), .B1(new_n766), .B2(new_n798), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n793), .B(new_n801), .C1(KEYINPUT92), .C2(new_n792), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n787), .B1(new_n790), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n756), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n759), .B1(new_n760), .B2(new_n803), .C1(new_n697), .C2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT93), .Z(new_n806));
  OAI21_X1  g0606(.A(new_n748), .B1(new_n697), .B2(G330), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n702), .B2(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n597), .A2(new_n692), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n606), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n668), .A2(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n682), .A2(new_n813), .A3(new_n692), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n813), .B(KEYINPUT98), .Z(new_n815));
  NAND2_X1  g0615(.A1(new_n682), .A2(new_n692), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n734), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n748), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n818), .B2(new_n819), .ZN(new_n823));
  INV_X1    g0623(.A(new_n813), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n754), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n760), .A2(new_n755), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n822), .B1(G77), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT94), .Z(new_n828));
  AOI22_X1  g0628(.A1(G283), .A2(new_n776), .B1(new_n780), .B2(G303), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n289), .B2(new_n781), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT95), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n763), .A2(new_n224), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G311), .B2(new_n767), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n283), .C1(new_n230), .C2(new_n770), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n795), .B(new_n834), .C1(G294), .C2(new_n773), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT96), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G137), .A2(new_n780), .B1(new_n776), .B2(G150), .ZN(new_n838));
  INV_X1    g0638(.A(G143), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n772), .C1(new_n798), .C2(new_n781), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n283), .B1(new_n791), .B2(G50), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n764), .A2(G68), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n766), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G58), .B2(new_n786), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n841), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n842), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n836), .A2(KEYINPUT96), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n837), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n828), .B1(new_n852), .B2(new_n757), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n821), .A2(new_n823), .B1(new_n825), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  NAND2_X1  g0655(.A1(new_n720), .A2(new_n733), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n676), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT101), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT40), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n579), .A2(new_n691), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n543), .A2(new_n584), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(new_n543), .B2(new_n584), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n813), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n720), .B2(new_n733), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n641), .A2(new_n634), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n295), .C1(new_n866), .C2(KEYINPUT16), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n641), .B2(new_n634), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT99), .B1(new_n868), .B2(new_n346), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n642), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n654), .ZN(new_n871));
  INV_X1    g0671(.A(new_n689), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n659), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n648), .A2(new_n653), .A3(new_n654), .ZN(new_n877));
  INV_X1    g0677(.A(new_n629), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n879), .B2(new_n873), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n655), .A2(new_n624), .A3(new_n628), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n655), .A2(new_n872), .ZN(new_n882));
  AND4_X1   g0682(.A1(new_n876), .A2(new_n881), .A3(new_n649), .A4(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n875), .B(KEYINPUT38), .C1(new_n880), .C2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n881), .A2(new_n882), .A3(new_n876), .A4(new_n649), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n649), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  INV_X1    g0687(.A(new_n882), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n885), .A2(new_n887), .B1(new_n659), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n884), .B1(KEYINPUT38), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n859), .B1(new_n864), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n871), .A2(new_n878), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n873), .A3(new_n649), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n883), .B1(new_n894), .B2(KEYINPUT37), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n659), .A2(new_n874), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT40), .B1(new_n897), .B2(new_n884), .ZN(new_n898));
  INV_X1    g0698(.A(new_n863), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n856), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n700), .B1(new_n858), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT102), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n902), .A2(new_n903), .B1(new_n858), .B2(new_n901), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n903), .B2(new_n902), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n890), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n584), .A2(new_n691), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n872), .B1(new_n644), .B2(new_n657), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n861), .A2(new_n862), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n668), .A2(new_n692), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n814), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n897), .A2(new_n884), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT100), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n911), .A2(new_n917), .A3(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n738), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n676), .B1(new_n923), .B2(new_n736), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n675), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n922), .B(new_n925), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n905), .A2(new_n926), .B1(new_n209), .B2(new_n742), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n905), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n426), .A2(new_n427), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(KEYINPUT35), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(G116), .A4(new_n220), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT36), .Z(new_n934));
  OAI211_X1 g0734(.A(new_n218), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n209), .B(G13), .C1(new_n935), .C2(new_n248), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n928), .A2(new_n934), .A3(new_n936), .ZN(G367));
  OR2_X1    g0737(.A1(new_n494), .A2(new_n692), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n497), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n490), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n449), .B(new_n451), .C1(new_n432), .C2(new_n692), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n433), .A2(new_n691), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n709), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT42), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n943), .A2(new_n368), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n691), .B1(new_n952), .B2(new_n449), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n946), .B2(KEYINPUT42), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n941), .B(new_n942), .C1(new_n951), .C2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n941), .A3(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT104), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n945), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n707), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n744), .B(KEYINPUT106), .ZN(new_n968));
  INV_X1    g0768(.A(new_n740), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n710), .A2(new_n945), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n710), .A2(new_n945), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT45), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(new_n707), .Z(new_n976));
  NAND3_X1  g0776(.A1(new_n699), .A2(new_n701), .A3(new_n705), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n707), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n685), .A3(new_n692), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n707), .A2(new_n708), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n969), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n713), .B(KEYINPUT41), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n968), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n967), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n750), .A2(new_n243), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n758), .C1(new_n213), .C2(new_n453), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n748), .B1(new_n987), .B2(KEYINPUT107), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(KEYINPUT107), .B2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(KEYINPUT46), .A2(G116), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n770), .A2(new_n990), .B1(new_n763), .B2(new_n292), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n280), .B(new_n991), .C1(G317), .C2(new_n767), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n770), .A2(new_n289), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(KEYINPUT46), .B2(new_n993), .C1(new_n230), .C2(new_n794), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT108), .B(G311), .Z(new_n995));
  AOI22_X1  g0795(.A1(G294), .A2(new_n776), .B1(new_n780), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G283), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n996), .B1(new_n997), .B2(new_n781), .C1(new_n281), .C2(new_n772), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G143), .A2(new_n780), .B1(new_n776), .B2(G159), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n201), .B2(new_n781), .C1(new_n558), .C2(new_n772), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n794), .A2(new_n203), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n283), .B1(new_n767), .B2(G137), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n791), .A2(G58), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n764), .A2(G77), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n994), .A2(new_n998), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n989), .B1(new_n1008), .B2(new_n757), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n804), .B2(new_n940), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n985), .A2(new_n1010), .ZN(G387));
  AOI21_X1  g0811(.A(new_n969), .B1(new_n979), .B2(new_n980), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n714), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n740), .B2(new_n981), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n968), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n981), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n213), .A2(new_n280), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n1017), .A2(new_n715), .B1(G107), .B2(new_n213), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n240), .A2(G45), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n750), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1021));
  NOR3_X1   g0821(.A1(new_n1021), .A2(G50), .A3(new_n557), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n260), .B1(new_n203), .B2(new_n228), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1022), .A2(G116), .A3(new_n462), .A4(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1021), .B1(G50), .B2(new_n557), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1018), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n758), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n822), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n283), .B1(new_n764), .B2(G97), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n791), .A2(G77), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n558), .C2(new_n766), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT110), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n794), .A2(new_n453), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n782), .B2(G68), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n776), .A2(new_n591), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G50), .A2(new_n773), .B1(new_n780), .B2(G159), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G322), .A2(new_n780), .B1(new_n776), .B2(new_n995), .ZN(new_n1039));
  INV_X1    g0839(.A(G317), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(new_n281), .B2(new_n781), .C1(new_n1040), .C2(new_n772), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(G294), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n794), .A2(new_n997), .B1(new_n770), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n280), .B1(new_n767), .B2(G326), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n289), .C2(new_n763), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT49), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1038), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1029), .B1(new_n1051), .B2(new_n757), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n706), .B2(new_n804), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1014), .A2(new_n1016), .A3(new_n1053), .ZN(G393));
  AOI21_X1  g0854(.A(new_n714), .B1(new_n976), .B2(new_n1012), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n976), .A2(new_n1012), .ZN(new_n1057));
  OAI21_X1  g0857(.A(KEYINPUT112), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT112), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1055), .B(new_n1059), .C1(new_n1012), .C2(new_n976), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n976), .A2(new_n1015), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n758), .B1(new_n292), .B2(new_n213), .C1(new_n1020), .C2(new_n247), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n822), .A2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n558), .A2(new_n779), .B1(new_n772), .B2(new_n798), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n794), .A2(new_n228), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n770), .A2(new_n203), .B1(new_n766), .B2(new_n839), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n283), .A4(new_n832), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n776), .B1(new_n782), .B2(new_n591), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1066), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G311), .A2(new_n773), .B1(new_n780), .B2(G317), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G283), .A2(new_n791), .B1(new_n767), .B2(G322), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n283), .A3(new_n797), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1044), .A2(new_n781), .B1(new_n775), .B2(new_n281), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n794), .A2(new_n289), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1071), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT111), .Z(new_n1080));
  OAI221_X1 g0880(.A(new_n1064), .B1(new_n804), .B2(new_n945), .C1(new_n1080), .C2(new_n760), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1061), .A2(new_n1062), .A3(new_n1081), .ZN(G390));
  AND3_X1   g0882(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n887), .A2(new_n885), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n660), .B2(new_n882), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n892), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n884), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1083), .A2(new_n1087), .B1(new_n915), .B2(new_n909), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n814), .A2(new_n914), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n908), .B(new_n890), .C1(new_n1090), .C2(new_n913), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n913), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n856), .A2(G330), .A3(new_n813), .A4(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n754), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n822), .B1(new_n591), .B2(new_n826), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n770), .A2(new_n558), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT53), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n794), .B2(new_n798), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1100), .B2(new_n1099), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT115), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1104), .A2(new_n782), .B1(new_n776), .B2(G137), .ZN(new_n1105));
  INV_X1    g0905(.A(G125), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n280), .B1(new_n766), .B2(new_n1106), .C1(new_n201), .C2(new_n763), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G132), .B2(new_n773), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n780), .A2(G128), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1102), .A2(new_n1105), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G107), .A2(new_n776), .B1(new_n780), .B2(G283), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n292), .B2(new_n781), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT116), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n844), .B1(new_n1044), .B2(new_n766), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n283), .B1(new_n770), .B2(new_n224), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1114), .A2(new_n1067), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(G116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n772), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1110), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1098), .B1(new_n1119), .B2(new_n757), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1096), .A2(new_n1015), .B1(new_n1097), .B2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT117), .Z(new_n1122));
  INV_X1    g0922(.A(KEYINPUT114), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n674), .B1(new_n739), .B2(new_n676), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT113), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n734), .A2(new_n676), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n700), .B(new_n664), .C1(new_n720), .C2(new_n733), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT113), .B1(new_n925), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n331), .A2(new_n376), .A3(new_n692), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n445), .A2(new_n452), .A3(new_n497), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT85), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n500), .A2(new_n377), .A3(new_n452), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n733), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n813), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1090), .B1(new_n1136), .B2(new_n913), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1092), .B1(new_n734), .B2(new_n815), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n913), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1090), .B1(new_n1140), .B2(new_n1093), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1127), .B(new_n1129), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1093), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1123), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n734), .A2(new_n815), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1090), .B(new_n1093), .C1(new_n1149), .C2(new_n1092), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1140), .A2(new_n1093), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1089), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n925), .A2(new_n1128), .A3(KEYINPUT113), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1125), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1096), .A2(new_n1153), .A3(new_n1156), .A4(KEYINPUT114), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1148), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1142), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n713), .C1(new_n1096), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1122), .A2(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1129), .A2(new_n1127), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT120), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1129), .A2(KEYINPUT120), .A3(new_n1127), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1148), .B2(new_n1157), .ZN(new_n1168));
  OAI21_X1  g0968(.A(G330), .B1(new_n891), .B2(new_n900), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n920), .A3(new_n921), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n890), .B(new_n899), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT40), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n864), .A2(new_n898), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n700), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n911), .A2(new_n917), .A3(KEYINPUT100), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT100), .B1(new_n911), .B2(new_n917), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n565), .A2(new_n689), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n578), .B(new_n1179), .Z(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(KEYINPUT119), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1178), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1170), .A2(new_n1177), .A3(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1162), .B1(new_n1168), .B2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1168), .A2(new_n1188), .A3(new_n1162), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n713), .B(new_n1189), .C1(new_n1190), .C2(KEYINPUT121), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1168), .A2(new_n1188), .A3(new_n1192), .A4(new_n1162), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1188), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1182), .A2(new_n754), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n822), .B1(G50), .B2(new_n826), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G58), .A2(new_n764), .B1(new_n767), .B2(G283), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n280), .A2(G41), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1031), .A3(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT118), .Z(new_n1201));
  OAI21_X1  g1001(.A(new_n1002), .B1(new_n292), .B2(new_n775), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G116), .A2(new_n780), .B1(new_n782), .B2(new_n454), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n230), .B2(new_n772), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G132), .A2(new_n776), .B1(new_n782), .B2(G137), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G125), .A2(new_n780), .B1(new_n773), .B2(G128), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1104), .A2(new_n791), .B1(G150), .B2(new_n786), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n270), .B(new_n504), .C1(new_n763), .C2(new_n798), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G124), .B2(new_n767), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1205), .A2(KEYINPUT58), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1199), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1218), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1206), .A2(new_n1216), .A3(new_n1217), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1197), .B1(new_n1220), .B2(new_n757), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1195), .A2(new_n1015), .B1(new_n1196), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1194), .A2(new_n1222), .ZN(G375));
  NAND3_X1  g1023(.A1(new_n1163), .A2(new_n1152), .A3(new_n1150), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n983), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1142), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n913), .A2(new_n754), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT122), .Z(new_n1228));
  OAI21_X1  g1028(.A(new_n822), .B1(G68), .B2(new_n826), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G283), .A2(new_n773), .B1(new_n780), .B2(G294), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n230), .B2(new_n781), .C1(new_n289), .C2(new_n775), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1034), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n791), .B1(new_n767), .B2(G303), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n283), .A3(new_n1005), .A4(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1104), .A2(new_n776), .B1(new_n773), .B2(G137), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n845), .B2(new_n779), .C1(new_n558), .C2(new_n781), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G159), .A2(new_n791), .B1(new_n767), .B2(G128), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n283), .B1(new_n764), .B2(G58), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n201), .C2(new_n794), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1231), .A2(new_n1234), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1229), .B1(new_n1240), .B2(new_n757), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1153), .A2(new_n1015), .B1(new_n1228), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1226), .A2(new_n1242), .ZN(G381));
  INV_X1    g1043(.A(G375), .ZN(new_n1244));
  OR3_X1    g1044(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G378), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n690), .A2(G213), .ZN(new_n1249));
  OR3_X1    g1049(.A1(G375), .A2(G378), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(G407), .A3(G213), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1250), .A2(G407), .A3(KEYINPUT123), .A4(G213), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G409));
  XNOR2_X1  g1055(.A(G393), .B(G396), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G390), .A2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n1061), .A3(new_n1062), .A4(new_n1081), .ZN(new_n1259));
  INV_X1    g1059(.A(G387), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1260), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1222), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1168), .A2(new_n1188), .A3(new_n983), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1222), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1247), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1224), .B1(new_n1159), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(KEYINPUT124), .B(new_n1224), .C1(new_n1159), .C2(new_n1272), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1224), .A2(new_n1272), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(new_n714), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1242), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n854), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(G384), .A3(new_n1242), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1270), .A2(new_n1271), .A3(new_n1249), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1266), .A2(new_n1269), .B1(G213), .B2(new_n690), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1283), .A2(G213), .A3(new_n690), .A4(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(G2897), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1281), .B(new_n1282), .C1(new_n1289), .C2(new_n1249), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1285), .B(new_n1286), .C1(new_n1287), .C2(new_n1291), .ZN(new_n1292));
  XOR2_X1   g1092(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(new_n1287), .B2(new_n1284), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1265), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1270), .A2(new_n1249), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1297), .B2(new_n1283), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1298), .A2(new_n1264), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1302), .ZN(G405));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1247), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1283), .A3(new_n1266), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G378), .B1(new_n1194), .B2(new_n1222), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1266), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1284), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1263), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(KEYINPUT126), .A3(new_n1261), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1309), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1264), .A2(new_n1305), .A3(KEYINPUT126), .A4(new_n1308), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(G402));
endmodule


