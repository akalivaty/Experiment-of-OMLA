//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n445, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(G217));
  NAND4_X1  g028(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n462), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n464), .A2(new_n466), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(G2105), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n462), .A3(new_n482), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n481), .A2(new_n490), .A3(new_n462), .A4(new_n482), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n492), .B2(G136), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n464), .A2(new_n466), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n465), .A2(G2104), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n462), .A2(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT4), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n467), .B2(new_n468), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n462), .B1(new_n499), .B2(new_n500), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n519), .ZN(G164));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n522), .A2(new_n523), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT5), .B(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G62), .ZN(new_n535));
  NAND2_X1  g110(.A1(G75), .A2(G543), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT73), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n532), .A2(new_n538), .ZN(G166));
  AOI22_X1  g114(.A1(new_n521), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n522), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n541), .A2(new_n534), .B1(new_n542), .B2(G51), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  AOI22_X1  g122(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n533), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n522), .A2(new_n550), .B1(new_n530), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n549), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND3_X1  g129(.A1(new_n521), .A2(G43), .A3(G543), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(new_n530), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n534), .A2(G56), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n533), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G188));
  NAND3_X1  g143(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT75), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n571), .B(KEYINPUT9), .C1(KEYINPUT75), .C2(new_n569), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n530), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n534), .A2(new_n521), .A3(KEYINPUT77), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G91), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  OAI211_X1 g153(.A(KEYINPUT75), .B(new_n578), .C1(new_n569), .C2(new_n570), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n534), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n533), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n572), .A2(new_n577), .A3(new_n579), .A4(new_n581), .ZN(G299));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n576), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n542), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NOR2_X1   g162(.A1(new_n530), .A2(new_n573), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT77), .B1(new_n534), .B2(new_n521), .ZN(new_n589));
  OAI21_X1  g164(.A(G86), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n576), .A2(new_n592), .A3(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n534), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n542), .B2(G48), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n594), .A2(new_n599), .ZN(G305));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT79), .B(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n522), .A2(new_n601), .B1(new_n530), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n533), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n576), .A2(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n534), .A2(G66), .ZN(new_n612));
  INV_X1    g187(.A(G79), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n613), .B2(new_n524), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n613), .A2(new_n524), .A3(KEYINPUT81), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(new_n542), .B2(G54), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n576), .A2(new_n618), .A3(G92), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n611), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n609), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n609), .B1(new_n621), .B2(G868), .ZN(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(G299), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n624), .B2(G168), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n624), .B2(G168), .ZN(G280));
  INV_X1    g202(.A(G860), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n620), .B1(G559), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT82), .ZN(G148));
  OR2_X1    g205(.A1(new_n620), .A2(G559), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n509), .A2(new_n474), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2100), .Z(new_n638));
  AND2_X1   g213(.A1(new_n492), .A2(G135), .ZN(new_n639));
  INV_X1    g214(.A(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n642));
  OAI22_X1  g217(.A1(new_n483), .A2(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n638), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2435), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2438), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n680), .A2(KEYINPUT83), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(KEYINPUT83), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n683), .A2(new_n684), .B1(new_n677), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n676), .A3(new_n680), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n688), .C1(new_n684), .C2(new_n683), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT84), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT85), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  AND2_X1   g273(.A1(KEYINPUT88), .A2(G16), .ZN(new_n699));
  NOR2_X1   g274(.A1(KEYINPUT88), .A2(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G6), .B(G305), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G16), .B2(G23), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n713), .A2(G1976), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(G1976), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n706), .B(new_n709), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n717), .B2(KEYINPUT34), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G25), .A2(G29), .ZN(new_n724));
  INV_X1    g299(.A(new_n483), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G119), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT86), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n492), .A2(G131), .ZN(new_n728));
  NOR2_X1   g303(.A1(G95), .A2(G2105), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT87), .Z(new_n732));
  AOI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT35), .B(G1991), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G24), .B(G290), .S(new_n701), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n723), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(KEYINPUT36), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n723), .A2(new_n742), .A3(new_n736), .A4(new_n739), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT94), .B1(new_n745), .B2(G29), .ZN(new_n746));
  OR3_X1    g321(.A1(new_n745), .A2(KEYINPUT94), .A3(G29), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n746), .B(new_n747), .C1(G162), .C2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT29), .Z(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(KEYINPUT95), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(KEYINPUT95), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n752), .B(new_n753), .Z(new_n754));
  OR2_X1    g329(.A1(G104), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n756));
  INV_X1    g331(.A(G128), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n483), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n492), .B2(G140), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n748), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n748), .A2(G26), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT28), .B2(new_n761), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G2067), .Z(new_n764));
  NAND2_X1  g339(.A1(G299), .A2(G16), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n767));
  INV_X1    g342(.A(G20), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n701), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G1956), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT30), .B(G28), .Z(new_n773));
  OAI211_X1 g348(.A(new_n764), .B(new_n772), .C1(G29), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n702), .A2(G19), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n561), .B2(new_n702), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1341), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n639), .A2(new_n748), .A3(new_n643), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G32), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT26), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n492), .B2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n474), .A2(G105), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n725), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT27), .B(G1996), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n492), .A2(G139), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n509), .A2(G127), .ZN(new_n791));
  AND2_X1   g366(.A1(G115), .A2(G2104), .ZN(new_n792));
  OAI21_X1  g367(.A(G2105), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  NAND3_X1  g370(.A1(new_n790), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G33), .B(new_n796), .S(G29), .Z(new_n797));
  OAI21_X1  g372(.A(new_n789), .B1(G2072), .B2(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n774), .A2(new_n777), .A3(new_n778), .A4(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G5), .B(G301), .S(G16), .Z(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT92), .Z(new_n801));
  INV_X1    g376(.A(G1961), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n621), .A2(G16), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G4), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G34), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(KEYINPUT24), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(KEYINPUT24), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n748), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G160), .B2(new_n748), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(G2084), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n799), .A2(new_n803), .A3(new_n807), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n797), .A2(G2072), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  INV_X1    g391(.A(G21), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G286), .B2(G16), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT91), .Z(new_n820));
  AOI22_X1  g395(.A1(new_n820), .A2(G1966), .B1(G2084), .B2(new_n812), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT31), .B(G11), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n805), .A2(new_n806), .ZN(new_n823));
  INV_X1    g398(.A(G27), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT93), .B1(new_n824), .B2(G29), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n824), .A2(KEYINPUT93), .A3(G29), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n826), .C1(G164), .C2(new_n748), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G2078), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(G2078), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n830), .B1(new_n820), .B2(G1966), .C1(new_n801), .C2(new_n802), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n814), .A2(new_n816), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n744), .A2(new_n754), .A3(new_n832), .ZN(G311));
  NAND3_X1  g408(.A1(new_n744), .A2(new_n754), .A3(new_n832), .ZN(G150));
  XNOR2_X1  g409(.A(KEYINPUT96), .B(G55), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n521), .A2(new_n835), .A3(G543), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n836), .B1(new_n837), .B2(new_n530), .C1(new_n838), .C2(new_n533), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT99), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n621), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n838), .A2(new_n533), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n836), .B1(new_n837), .B2(new_n530), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n555), .B1(new_n556), .B2(new_n530), .C1(new_n850), .C2(new_n533), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n846), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n839), .A2(new_n561), .A3(KEYINPUT97), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n839), .B2(new_n561), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n849), .A2(new_n851), .A3(KEYINPUT98), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n845), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n842), .B1(new_n860), .B2(G860), .ZN(G145));
  XOR2_X1   g436(.A(new_n644), .B(G160), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n796), .B(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n636), .ZN(new_n867));
  INV_X1    g442(.A(new_n759), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n492), .A2(new_n869), .A3(G142), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n492), .B2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  INV_X1    g449(.A(G118), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n463), .B1(new_n875), .B2(G2105), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n725), .A2(G130), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n868), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n492), .A2(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n877), .A3(new_n870), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(new_n759), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n785), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n873), .A2(new_n868), .A3(new_n877), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n759), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n786), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n883), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n867), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n887), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n786), .B1(new_n885), .B2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT102), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n636), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n515), .A2(new_n517), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n731), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n890), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n890), .B2(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n866), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n888), .A2(new_n889), .A3(new_n867), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n636), .B1(new_n893), .B2(new_n894), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n897), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n863), .B(new_n864), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n890), .A2(new_n895), .A3(new_n898), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g485(.A1(new_n839), .A2(G868), .ZN(new_n911));
  NOR2_X1   g486(.A1(G299), .A2(new_n620), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n620), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(G299), .A2(new_n620), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT41), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT103), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n920), .B(KEYINPUT41), .C1(new_n917), .C2(new_n912), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n859), .B(new_n631), .Z(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n917), .A2(new_n912), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G288), .B(G303), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(G290), .ZN(new_n931));
  INV_X1    g506(.A(G305), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n924), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n931), .B(G305), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n928), .A3(new_n927), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n911), .B1(new_n940), .B2(G868), .ZN(G295));
  XOR2_X1   g516(.A(G295), .B(KEYINPUT105), .Z(G331));
  AND3_X1   g517(.A1(new_n854), .A2(new_n858), .A3(G301), .ZN(new_n943));
  AOI21_X1  g518(.A(G301), .B1(new_n854), .B2(new_n858), .ZN(new_n944));
  OAI21_X1  g519(.A(G286), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n859), .A2(G171), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n854), .A2(new_n858), .A3(G301), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(G168), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n948), .A3(new_n925), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT107), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n945), .A2(new_n948), .A3(new_n951), .A4(new_n925), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n945), .A2(new_n948), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n956), .B2(new_n922), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n955), .A2(KEYINPUT106), .A3(new_n921), .A4(new_n919), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n937), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n945), .A2(new_n948), .B1(new_n918), .B2(new_n916), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n949), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n933), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n957), .A2(new_n958), .ZN(new_n967));
  INV_X1    g542(.A(new_n953), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n933), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT43), .B1(new_n960), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT44), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n960), .B2(new_n970), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n967), .A2(new_n968), .A3(new_n937), .ZN(new_n975));
  AND4_X1   g550(.A1(new_n973), .A2(new_n975), .A3(new_n902), .A4(new_n965), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(KEYINPUT44), .B2(new_n977), .ZN(G397));
  NOR2_X1   g553(.A1(new_n479), .A2(G2105), .ZN(new_n979));
  AOI22_X1  g554(.A1(G101), .A2(new_n474), .B1(new_n979), .B2(G137), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n509), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n981));
  OAI211_X1 g556(.A(G40), .B(new_n980), .C1(new_n981), .C2(new_n462), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n515), .B2(new_n517), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT45), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n731), .B(new_n734), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n785), .B(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n759), .B(G2067), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NOR2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n592), .B1(new_n576), .B2(G86), .ZN(new_n997));
  INV_X1    g572(.A(G86), .ZN(new_n998));
  AOI211_X1 g573(.A(KEYINPUT78), .B(new_n998), .C1(new_n574), .C2(new_n575), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n996), .B(new_n599), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT114), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n594), .A2(new_n1002), .A3(new_n996), .A4(new_n599), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n534), .A2(new_n521), .A3(G86), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n996), .B1(new_n599), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(G8), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n896), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(new_n982), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G40), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n471), .A2(new_n477), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n983), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(KEYINPUT113), .A3(new_n1011), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1004), .A2(KEYINPUT49), .A3(new_n1007), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1010), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n710), .A2(G1976), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n1031));
  OAI21_X1  g606(.A(G8), .B1(new_n532), .B2(new_n538), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(KEYINPUT110), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(G8), .C1(new_n532), .C2(new_n538), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(KEYINPUT110), .A3(new_n1031), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1035), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1038), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1033), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n1044));
  AOI211_X1 g619(.A(new_n1044), .B(G1384), .C1(new_n515), .C2(new_n517), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n512), .A2(new_n1012), .A3(new_n519), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n982), .B(new_n1045), .C1(new_n1046), .C2(new_n1044), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n982), .B1(new_n983), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1047), .A2(G1971), .B1(new_n1052), .B2(G2090), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n1053), .B2(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n995), .B1(new_n1030), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT49), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1009), .B(new_n1006), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1058), .A2(new_n1021), .B1(KEYINPUT52), .B2(new_n1025), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n982), .B1(new_n1046), .B2(new_n1044), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1045), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1971), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1048), .A2(new_n751), .A3(new_n1051), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1043), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1059), .A2(KEYINPUT117), .A3(new_n1029), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n896), .A2(new_n1012), .A3(new_n1050), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1018), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(KEYINPUT50), .B2(new_n1046), .ZN(new_n1070));
  INV_X1    g645(.A(G2084), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n982), .B1(new_n1013), .B2(new_n1044), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n1012), .A4(new_n519), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1070), .A2(new_n1071), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1011), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1076), .A2(G286), .A3(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1055), .A2(new_n1067), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1043), .B(G8), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n982), .B1(new_n1013), .B2(new_n1049), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n512), .A2(new_n1085), .A3(new_n1012), .A4(new_n519), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n751), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1047), .B2(G1971), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT116), .B(new_n1043), .C1(new_n1088), .C2(new_n1011), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1087), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1011), .B1(new_n1062), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1092), .B2(new_n1065), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1080), .A2(new_n1023), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1096), .A3(new_n1078), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1079), .A2(new_n1083), .B1(new_n1082), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1046), .A2(new_n1044), .ZN(new_n1099));
  INV_X1    g674(.A(G2078), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(new_n1061), .A3(new_n1100), .A4(new_n1018), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1052), .A2(new_n802), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1072), .A2(KEYINPUT53), .A3(new_n1100), .A4(new_n1073), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G171), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G168), .A2(new_n1077), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1108), .B(new_n1110), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1111));
  INV_X1    g686(.A(G8), .ZN(new_n1112));
  AND4_X1   g687(.A1(KEYINPUT45), .A2(new_n512), .A3(new_n1012), .A4(new_n519), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1018), .B1(KEYINPUT45), .B2(new_n983), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1075), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1048), .A2(new_n1071), .A3(new_n1051), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT51), .B1(new_n1117), .B2(new_n1109), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1076), .A2(new_n1110), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1111), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1107), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1095), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1111), .B(KEYINPUT62), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1059), .A2(new_n1081), .A3(new_n1029), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1023), .A2(new_n1027), .A3(new_n710), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1004), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(KEYINPUT115), .A3(new_n1004), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(new_n1021), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1125), .A2(new_n1126), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1098), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1047), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(G299), .B(KEYINPUT57), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(new_n771), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT118), .B(G1956), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1136), .B(new_n1138), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1136), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1144), .A2(KEYINPUT119), .A3(new_n1137), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT119), .B1(new_n1144), .B2(new_n1137), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1019), .A2(G2067), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1052), .B2(new_n806), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(new_n620), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1143), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  AOI21_X1  g727(.A(G1956), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(new_n1139), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1138), .B1(new_n1154), .B2(new_n1136), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1143), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT120), .B(new_n1152), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1143), .A2(KEYINPUT61), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n620), .B(KEYINPUT121), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1149), .A2(KEYINPUT60), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1149), .A2(KEYINPUT60), .B1(KEYINPUT121), .B2(new_n621), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT58), .B(G1341), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1019), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(G1996), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n561), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT59), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1163), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1151), .B1(new_n1161), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1103), .A2(G301), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT54), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1101), .A2(new_n1102), .B1(new_n1052), .B2(new_n802), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1072), .A2(KEYINPUT53), .A3(new_n1100), .A4(new_n1061), .ZN(new_n1181));
  AOI21_X1  g756(.A(G301), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(new_n1120), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1180), .A2(G301), .A3(new_n1181), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT54), .B1(new_n1107), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1186), .A2(KEYINPUT122), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1188), .B(KEYINPUT54), .C1(new_n1107), .C2(new_n1185), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1184), .B(new_n1123), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n994), .B1(new_n1134), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n984), .A2(new_n986), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT46), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n988), .A2(new_n786), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n984), .B2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT124), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT47), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n989), .A2(new_n984), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1201), .A2(new_n732), .A3(new_n735), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(G2067), .B2(new_n868), .ZN(new_n1203));
  OR2_X1    g778(.A1(new_n1203), .A2(KEYINPUT123), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(KEYINPUT123), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1204), .A2(new_n984), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n992), .A2(new_n984), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT48), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n990), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1200), .A2(new_n1206), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT125), .B1(new_n1193), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n994), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1097), .A2(new_n1082), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1055), .A2(new_n1067), .A3(new_n1078), .A4(new_n1083), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1215), .A2(new_n1126), .A3(new_n1132), .A4(new_n1125), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1144), .A2(new_n1137), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT119), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1144), .A2(KEYINPUT119), .A3(new_n1137), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1168), .B1(new_n1221), .B2(new_n1162), .ZN(new_n1222));
  NAND4_X1  g797(.A1(new_n1222), .A2(new_n1175), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1190), .B1(new_n1223), .B2(new_n1151), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1212), .B1(new_n1216), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1226));
  INV_X1    g801(.A(new_n1210), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1211), .A2(new_n1228), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1231));
  OAI21_X1  g805(.A(new_n697), .B1(new_n974), .B2(new_n976), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n660), .A2(G319), .A3(new_n673), .ZN(new_n1233));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g809(.A1(new_n660), .A2(KEYINPUT126), .A3(G319), .A4(new_n673), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g811(.A1(new_n909), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g812(.A(new_n1231), .B1(new_n1232), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g813(.A1(new_n975), .A2(new_n902), .ZN(new_n1240));
  NOR2_X1   g814(.A1(new_n959), .A2(new_n937), .ZN(new_n1241));
  OAI21_X1  g815(.A(KEYINPUT43), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g816(.A1(new_n960), .A2(new_n973), .A3(new_n965), .ZN(new_n1243));
  AOI21_X1  g817(.A(G229), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g818(.A1(new_n1244), .A2(KEYINPUT127), .A3(new_n909), .A4(new_n1237), .ZN(new_n1245));
  AND2_X1   g819(.A1(new_n1239), .A2(new_n1245), .ZN(G308));
  NAND2_X1  g820(.A1(new_n1239), .A2(new_n1245), .ZN(G225));
endmodule


