//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988;
  AND2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G169gat), .B2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT24), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n204), .A2(new_n210), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n204), .A2(new_n210), .A3(new_n215), .A4(KEYINPUT25), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G113gat), .B(G120gat), .Z(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g021(.A(G127gat), .B(G134gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n222), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(G134gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G127gat), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n225), .A2(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT26), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n214), .B(new_n233), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n237), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n241), .B(KEYINPUT65), .C1(new_n237), .C2(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT64), .B(KEYINPUT28), .C1(new_n246), .C2(G190gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n243), .A4(new_n245), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n240), .A2(new_n242), .A3(new_n247), .A4(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n232), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n232), .B1(new_n220), .B2(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(G227gat), .ZN(new_n256));
  INV_X1    g055(.A(G233gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n258), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n220), .A2(new_n252), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n224), .A2(new_n231), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n266), .B1(new_n269), .B2(new_n253), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT32), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT67), .B1(new_n270), .B2(KEYINPUT33), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n258), .B1(new_n254), .B2(new_n255), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT33), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n265), .A2(KEYINPUT33), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n261), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n264), .B1(new_n274), .B2(KEYINPUT32), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n270), .A2(KEYINPUT67), .A3(KEYINPUT33), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(new_n280), .A3(new_n260), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n259), .B2(KEYINPUT68), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n282), .B2(new_n287), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G211gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT70), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G211gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT22), .B1(new_n300), .B2(G218gat), .ZN(new_n301));
  XOR2_X1   g100(.A(G197gat), .B(G204gat), .Z(new_n302));
  OAI21_X1  g101(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT70), .B(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n302), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n294), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G141gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n320), .A3(G148gat), .ZN(new_n321));
  INV_X1    g120(.A(G148gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G141gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(G162gat), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT2), .B1(new_n325), .B2(new_n314), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n317), .A2(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n316), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n327), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n311), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G228gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n257), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n324), .A2(new_n326), .B1(new_n316), .B2(new_n331), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT3), .B1(new_n310), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n337), .B(new_n339), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n294), .B1(new_n307), .B2(new_n308), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n336), .B1(new_n344), .B2(KEYINPUT82), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n303), .A2(new_n346), .A3(new_n309), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n333), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n337), .B1(new_n348), .B2(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350));
  INV_X1    g149(.A(new_n339), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n343), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n293), .B1(new_n354), .B2(G22gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G22gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n334), .ZN(new_n361));
  INV_X1    g160(.A(new_n336), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n310), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n303), .A2(new_n346), .A3(new_n309), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n303), .B2(new_n346), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n334), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n327), .A2(new_n332), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT83), .B1(new_n368), .B2(new_n339), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n360), .B1(new_n371), .B2(new_n343), .ZN(new_n372));
  INV_X1    g171(.A(new_n343), .ZN(new_n373));
  AOI211_X1 g172(.A(G22gat), .B(new_n373), .C1(new_n369), .C2(new_n370), .ZN(new_n374));
  OAI22_X1  g173(.A1(new_n355), .A2(new_n359), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n354), .A2(G22gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n360), .A3(new_n343), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n293), .A4(new_n358), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n292), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n232), .B1(new_n367), .B2(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n361), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT78), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT4), .B1(new_n367), .B2(new_n268), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n340), .A2(new_n232), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n340), .A2(new_n232), .A3(KEYINPUT81), .A4(new_n391), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n340), .A2(new_n232), .A3(new_n397), .A4(new_n391), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n385), .B1(new_n381), .B2(new_n361), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n340), .B(new_n232), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n383), .B1(new_n402), .B2(new_n385), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n388), .A2(new_n395), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(G1gat), .B(G29gat), .Z(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT86), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT6), .B1(new_n404), .B2(new_n409), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n401), .A2(new_n403), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n400), .A2(new_n393), .A3(new_n383), .A4(new_n394), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(KEYINPUT6), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT35), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G8gat), .B(G36gat), .Z(new_n420));
  XOR2_X1   g219(.A(G64gat), .B(G92gat), .Z(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n267), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n220), .A2(KEYINPUT72), .A3(new_n252), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n267), .A2(new_n425), .A3(new_n362), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n311), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n267), .A2(new_n425), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n427), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n426), .A2(KEYINPUT29), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n422), .B(new_n430), .C1(new_n434), .C2(new_n311), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n433), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n424), .B2(new_n427), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n310), .B1(new_n439), .B2(new_n431), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n422), .A4(new_n430), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n430), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n422), .B(KEYINPUT73), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n437), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n437), .A2(new_n444), .A3(KEYINPUT85), .A4(new_n441), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n419), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n412), .A2(new_n409), .A3(new_n413), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n418), .B1(new_n453), .B2(new_n414), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n437), .A2(new_n444), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n441), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n292), .A2(new_n379), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n380), .A2(new_n450), .B1(new_n458), .B2(KEYINPUT35), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n462), .C1(new_n290), .C2(new_n291), .ZN(new_n463));
  INV_X1    g262(.A(new_n289), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n278), .A2(new_n281), .A3(new_n261), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n260), .B1(new_n286), .B2(new_n280), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(KEYINPUT69), .A3(new_n460), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n456), .A2(new_n375), .A3(new_n378), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n414), .A2(new_n415), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT86), .B(new_n409), .C1(new_n412), .C2(new_n413), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT39), .B1(new_n402), .B2(new_n385), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n393), .A2(new_n382), .A3(new_n394), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n385), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n480), .A3(new_n385), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n409), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n409), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT40), .B1(new_n483), .B2(new_n477), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n447), .A2(new_n448), .A3(new_n474), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n440), .A2(new_n487), .A3(new_n430), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n428), .A2(new_n310), .A3(new_n429), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(KEYINPUT37), .C1(new_n434), .C2(new_n310), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n443), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(new_n435), .ZN(new_n494));
  INV_X1    g293(.A(new_n422), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n487), .B1(new_n440), .B2(new_n430), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT38), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n417), .A3(new_n418), .A4(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n379), .A2(new_n486), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n471), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT87), .B1(new_n459), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n450), .A2(new_n379), .A3(new_n292), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n379), .A2(new_n486), .A3(new_n499), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n507), .A2(new_n470), .A3(new_n469), .A4(new_n463), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(G1gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(G1gat), .B2(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  INV_X1    g319(.A(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT14), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT88), .B1(new_n523), .B2(new_n525), .ZN(new_n529));
  OAI211_X1 g328(.A(KEYINPUT15), .B(new_n519), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT89), .B(G50gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(G43gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n534));
  INV_X1    g333(.A(new_n526), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n520), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n530), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n538), .A2(new_n542), .A3(new_n540), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n530), .A2(KEYINPUT17), .A3(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n517), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n511), .B(new_n541), .C1(new_n543), .C2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT18), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT12), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n546), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n511), .B(KEYINPUT13), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n540), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n517), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n560), .B2(new_n541), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n549), .A2(new_n554), .A3(new_n556), .A4(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n561), .B1(new_n548), .B2(KEYINPUT18), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n554), .B1(new_n565), .B2(new_n556), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n575));
  INV_X1    g374(.A(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G99gat), .ZN(new_n579));
  INV_X1    g378(.A(G106gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT8), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT7), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n574), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n578), .A3(new_n581), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(new_n573), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n572), .B1(new_n559), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n544), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n543), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n570), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n543), .A2(new_n592), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n599), .B2(new_n590), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(new_n569), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n598), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n598), .B2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n611));
  OR2_X1    g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G64gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G57gat), .ZN(new_n617));
  INV_X1    g416(.A(G57gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G64gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(KEYINPUT92), .B2(KEYINPUT9), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT9), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n610), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n618), .B2(G64gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n616), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n626), .A3(new_n619), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n615), .A2(new_n621), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G127gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n621), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n623), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT95), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(KEYINPUT21), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n517), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n632), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT94), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G155gat), .ZN(new_n644));
  XOR2_X1   g443(.A(G183gat), .B(G211gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n641), .B(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n635), .B1(new_n585), .B2(new_n587), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n582), .A2(new_n574), .A3(new_n584), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n586), .A2(new_n573), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n628), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n588), .A2(new_n636), .A3(KEYINPUT10), .A4(new_n638), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G230gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n257), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  AND2_X1   g461(.A1(new_n648), .A2(new_n652), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n659), .B(new_n662), .C1(new_n658), .C2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n662), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n657), .B1(new_n653), .B2(new_n654), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n663), .A2(new_n658), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n609), .A2(new_n647), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n510), .A2(new_n568), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT98), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n510), .A2(new_n675), .A3(new_n568), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n454), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  INV_X1    g479(.A(new_n449), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND4_X1   g481(.A1(KEYINPUT42), .A2(new_n677), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n677), .B2(new_n681), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT99), .B(new_n449), .C1(new_n674), .C2(new_n676), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(G8gat), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT100), .A4(new_n516), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n677), .A2(new_n695), .A3(new_n292), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n463), .A2(new_n469), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n674), .B2(new_n676), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n699), .B2(new_n695), .ZN(G1326gat));
  INV_X1    g499(.A(new_n379), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n677), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n609), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n459), .A2(new_n501), .A3(KEYINPUT87), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n506), .B1(new_n505), .B2(new_n508), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n505), .A2(new_n508), .ZN(new_n710));
  INV_X1    g509(.A(new_n608), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n606), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n705), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n564), .B2(new_n566), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n549), .A2(new_n556), .A3(new_n562), .ZN(new_n719));
  INV_X1    g518(.A(new_n554), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(KEYINPUT102), .A3(new_n563), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n647), .A2(new_n669), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n716), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n454), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n712), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT101), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n510), .A2(new_n568), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n521), .A3(new_n678), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n728), .A2(new_n734), .A3(new_n735), .ZN(G1328gat));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n522), .A3(new_n681), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n737), .B(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G36gat), .B1(new_n727), .B2(new_n449), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n740), .B(new_n741), .C1(new_n738), .C2(KEYINPUT46), .ZN(G1329gat));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n731), .A2(new_n743), .A3(new_n292), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n709), .A2(new_n697), .A3(new_n714), .A4(new_n726), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G43gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n744), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT105), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n744), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n747), .B(new_n754), .ZN(G1330gat));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n532), .B1(new_n727), .B2(new_n379), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n379), .A2(new_n532), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n731), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1331gat));
  NAND3_X1  g564(.A1(new_n609), .A2(new_n647), .A3(new_n669), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n723), .B(new_n766), .C1(new_n505), .C2(new_n508), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n678), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g568(.A(new_n449), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n772), .B(new_n773), .Z(G1333gat));
  AND2_X1   g573(.A1(new_n767), .A2(new_n292), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(KEYINPUT109), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(KEYINPUT109), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n776), .A2(new_n777), .A3(G71gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n767), .A2(G71gat), .A3(new_n697), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n767), .A2(new_n701), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n575), .A2(new_n577), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n723), .A2(new_n647), .A3(new_n670), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n715), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n788), .B2(new_n454), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n723), .A2(new_n647), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n712), .B(new_n791), .C1(new_n459), .C2(new_n501), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n609), .B1(new_n505), .B2(new_n508), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n791), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n794), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n792), .A2(new_n793), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n454), .A2(new_n784), .A3(new_n670), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n789), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n449), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n576), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n449), .A2(G92gat), .A3(new_n670), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n794), .A2(new_n797), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n800), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n802), .A2(new_n808), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n805), .B2(new_n576), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n788), .B2(new_n698), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n292), .A2(new_n579), .A3(new_n669), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n802), .B2(new_n817), .ZN(G1338gat));
  NAND4_X1  g617(.A1(new_n709), .A2(new_n701), .A3(new_n714), .A4(new_n785), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G106gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n701), .A2(new_n580), .A3(new_n669), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n809), .B2(new_n800), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(KEYINPUT112), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n824), .B(new_n821), .C1(new_n809), .C2(new_n800), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n820), .C1(new_n802), .C2(new_n821), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1339gat));
  NOR2_X1   g632(.A1(new_n723), .A2(new_n671), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n659), .A2(KEYINPUT54), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n662), .B1(new_n666), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n664), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n839), .A3(KEYINPUT55), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(new_n837), .B2(new_n839), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n664), .A3(new_n840), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(KEYINPUT115), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n543), .A2(new_n545), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n511), .B1(new_n850), .B2(new_n541), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n560), .A2(new_n541), .A3(new_n558), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n553), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n563), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n712), .A2(new_n846), .A3(new_n849), .A4(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n563), .A2(new_n669), .A3(new_n853), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT116), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n718), .A2(new_n722), .A3(new_n849), .A4(new_n846), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n609), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n835), .B1(new_n861), .B2(new_n647), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n380), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n681), .A2(new_n454), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n567), .ZN(new_n866));
  INV_X1    g665(.A(G113gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n723), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT117), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n865), .B2(new_n869), .ZN(G1340gat));
  NOR2_X1   g669(.A1(new_n865), .A2(new_n670), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(G120gat), .Z(G1341gat));
  INV_X1    g671(.A(new_n647), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g673(.A(KEYINPUT118), .B(G127gat), .Z(new_n875));
  XNOR2_X1  g674(.A(new_n874), .B(new_n875), .ZN(G1342gat));
  NOR2_X1   g675(.A1(new_n609), .A2(new_n681), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n863), .A2(new_n229), .A3(new_n678), .A4(new_n877), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT56), .Z(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n865), .B2(new_n609), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n318), .A2(new_n320), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n860), .A2(new_n609), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n647), .B1(new_n884), .B2(new_n855), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n883), .B(new_n701), .C1(new_n885), .C2(new_n834), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n698), .A2(new_n864), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n837), .A2(new_n839), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT119), .B1(new_n888), .B2(KEYINPUT55), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n847), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n889), .A2(new_n841), .A3(new_n845), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n857), .B1(new_n567), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n609), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n647), .B1(new_n894), .B2(new_n855), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n701), .B1(new_n895), .B2(new_n834), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n887), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n882), .B1(new_n898), .B2(new_n567), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(new_n887), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n567), .A2(G141gat), .ZN(new_n902));
  AND4_X1   g701(.A1(new_n701), .A2(new_n862), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n897), .A3(new_n723), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n882), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n904), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n909), .B2(KEYINPUT58), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n903), .B1(new_n907), .B2(new_n882), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(KEYINPUT120), .A3(new_n900), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n905), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT121), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n905), .C1(new_n910), .C2(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1344gat));
  AND2_X1   g716(.A1(new_n862), .A2(new_n701), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n901), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n322), .A3(new_n669), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n918), .A2(new_n883), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n671), .A2(new_n568), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n883), .B(new_n701), .C1(new_n895), .C2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n669), .A3(new_n901), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n898), .A2(new_n670), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(KEYINPUT59), .A3(new_n322), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n920), .B1(new_n927), .B2(new_n929), .ZN(G1345gat));
  NAND3_X1  g729(.A1(new_n919), .A2(new_n314), .A3(new_n647), .ZN(new_n931));
  OAI21_X1  g730(.A(G155gat), .B1(new_n898), .B2(new_n873), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1346gat));
  NAND2_X1  g732(.A1(new_n678), .A2(new_n325), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n698), .A3(new_n877), .A4(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n898), .A2(new_n609), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n325), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n449), .A2(new_n678), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n380), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n862), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n206), .A3(new_n723), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT122), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n206), .B1(new_n941), .B2(new_n568), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(G1348gat));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n669), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g746(.A1(new_n941), .A2(new_n647), .ZN(new_n948));
  MUX2_X1   g747(.A(new_n246), .B(new_n211), .S(new_n948), .Z(new_n949));
  XNOR2_X1  g748(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n949), .B(new_n950), .ZN(G1350gat));
  NAND2_X1  g750(.A1(new_n941), .A2(new_n712), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(G190gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(G190gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT125), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n955), .A2(KEYINPUT125), .A3(new_n957), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G1351gat));
  NAND2_X1  g762(.A1(new_n698), .A2(new_n939), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n918), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  AOI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n723), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n922), .A2(new_n924), .A3(new_n965), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(new_n567), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n968), .A2(new_n971), .ZN(G1352gat));
  NOR3_X1   g771(.A1(new_n966), .A2(G204gat), .A3(new_n670), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n969), .B2(new_n670), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n967), .A2(new_n305), .A3(new_n647), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n925), .A2(new_n647), .A3(new_n965), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n979));
  OAI211_X1 g778(.A(KEYINPUT63), .B(G211gat), .C1(new_n969), .C2(new_n873), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n977), .B1(new_n979), .B2(new_n981), .ZN(G1354gat));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n306), .A3(new_n712), .ZN(new_n983));
  OAI21_X1  g782(.A(G218gat), .B1(new_n969), .B2(new_n609), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n983), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(G1355gat));
endmodule


