//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n637,
    new_n640, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT64), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI21_X1  g031(.A(KEYINPUT65), .B1(new_n451), .B2(G2106), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n451), .A2(KEYINPUT65), .A3(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT3), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT67), .B1(new_n467), .B2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(new_n466), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OR3_X1    g047(.A1(new_n471), .A2(KEYINPUT68), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT68), .B1(new_n471), .B2(new_n472), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n464), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(new_n466), .A3(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n481), .A2(G2105), .B1(new_n484), .B2(G101), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n473), .A2(new_n474), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  OR3_X1    g063(.A1(new_n488), .A2(G100), .A3(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(G100), .B2(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n466), .A2(G112), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n489), .A2(new_n490), .A3(G2104), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G136), .ZN(new_n493));
  INV_X1    g068(.A(new_n470), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(new_n468), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(G2105), .A3(new_n465), .ZN(new_n496));
  INV_X1    g071(.A(G124), .ZN(new_n497));
  OAI221_X1 g072(.A(new_n492), .B1(new_n471), .B2(new_n493), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  INV_X1    g075(.A(new_n471), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G136), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(new_n492), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(G162));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR4_X1   g081(.A1(new_n479), .A2(KEYINPUT4), .A3(new_n506), .A4(G2105), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n495), .A2(G138), .A3(new_n465), .A4(new_n466), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n495), .A2(G126), .A3(new_n465), .A4(G2105), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n466), .A2(G114), .ZN(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  OR3_X1    g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT71), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT71), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(new_n516), .ZN(G164));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n519), .B2(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n520), .A2(new_n523), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n528), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n527), .B(new_n531), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT73), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n533), .A2(new_n528), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G88), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n538), .A2(new_n539), .A3(new_n527), .A4(new_n531), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(G166));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n530), .A2(G51), .B1(new_n533), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n528), .A2(G89), .A3(new_n520), .A4(new_n523), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n545), .B1(new_n544), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n543), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n543), .B(KEYINPUT75), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(G168));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n524), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n528), .A2(G90), .A3(new_n520), .A4(new_n523), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n528), .A2(G52), .A3(G543), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n559), .A2(KEYINPUT76), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT76), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  INV_X1    g139(.A(G81), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n534), .A2(new_n565), .B1(new_n566), .B2(new_n529), .ZN(new_n567));
  INV_X1    g142(.A(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n533), .A2(G56), .ZN(new_n569));
  NAND2_X1  g144(.A1(G68), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  AND3_X1   g148(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G36), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT77), .ZN(G188));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n529), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n537), .A2(G91), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT78), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT78), .B1(new_n520), .B2(new_n523), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n583), .B(new_n584), .C1(new_n568), .C2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G168), .ZN(G286));
  INV_X1    g165(.A(G166), .ZN(G303));
  NAND2_X1  g166(.A1(new_n530), .A2(G49), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n534), .ZN(G288));
  NAND2_X1  g170(.A1(new_n533), .A2(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n568), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n533), .A2(G86), .A3(new_n528), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n528), .A2(G48), .A3(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n537), .A2(G85), .B1(G47), .B2(new_n530), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n524), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n609), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n530), .A2(G54), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n587), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n617));
  OAI211_X1 g192(.A(KEYINPUT80), .B(new_n616), .C1(new_n617), .C2(new_n568), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n524), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT78), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(G66), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n568), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n616), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n537), .A2(G92), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT10), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n615), .B1(new_n632), .B2(G868), .ZN(G284));
  OAI21_X1  g208(.A(new_n615), .B1(new_n632), .B2(G868), .ZN(G321));
  NAND2_X1  g209(.A1(G286), .A2(G868), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(G868), .B2(new_n636), .ZN(new_n637));
  MUX2_X1   g212(.A(new_n635), .B(new_n637), .S(KEYINPUT81), .Z(G297));
  MUX2_X1   g213(.A(new_n635), .B(new_n637), .S(KEYINPUT81), .Z(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n632), .B1(new_n640), .B2(G860), .ZN(G148));
  OAI21_X1  g216(.A(G868), .B1(new_n631), .B2(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(G868), .B2(new_n572), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  INV_X1    g222(.A(G123), .ZN(new_n648));
  OAI221_X1 g223(.A(new_n646), .B1(new_n471), .B2(new_n647), .C1(new_n496), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT82), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  OR3_X1    g226(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n479), .ZN(new_n652));
  OAI21_X1  g227(.A(KEYINPUT12), .B1(new_n483), .B2(new_n479), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT13), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n656), .ZN(G156));
  XOR2_X1   g232(.A(KEYINPUT15), .B(G2435), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT83), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n663), .A3(KEYINPUT14), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT16), .B(G1341), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1348), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(G14), .B1(new_n664), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(G401));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  XNOR2_X1  g248(.A(G2084), .B(G2090), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n679), .A2(KEYINPUT17), .A3(new_n676), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n676), .B1(new_n679), .B2(KEYINPUT17), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n680), .A2(new_n681), .A3(new_n675), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT20), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n688), .A2(new_n692), .A3(new_n696), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n694), .A2(new_n695), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n703), .B(new_n706), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  NOR2_X1   g283(.A1(G16), .A2(G22), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G166), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1971), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G6), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n602), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G23), .B(G288), .S(G16), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n711), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT34), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n495), .A2(G119), .A3(new_n465), .A4(G2105), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n495), .A2(G131), .A3(new_n465), .A4(new_n466), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n466), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n724), .B2(new_n725), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n722), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(KEYINPUT89), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n722), .A2(new_n723), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT87), .B(G29), .ZN(new_n735));
  MUX2_X1   g310(.A(G25), .B(new_n734), .S(new_n735), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n736), .B(new_n737), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n712), .A2(G24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n613), .B2(new_n712), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1986), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n721), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n712), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n572), .B2(new_n712), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G1341), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G1341), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT30), .B(G28), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n754), .A2(G2072), .B1(G29), .B2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  INV_X1    g331(.A(G127), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n479), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2105), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n761), .C1(new_n471), .C2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n754), .A2(G2072), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n649), .B(KEYINPUT82), .ZN(new_n768));
  INV_X1    g343(.A(new_n735), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT27), .B(G1996), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n749), .A2(G32), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT26), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n484), .B2(G105), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n495), .A2(G141), .A3(new_n465), .A4(new_n466), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n495), .A2(G129), .A3(new_n465), .A4(G2105), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n772), .B1(new_n782), .B2(new_n749), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n753), .B(new_n770), .C1(new_n771), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n769), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n769), .ZN(new_n786));
  MUX2_X1   g361(.A(new_n785), .B(new_n786), .S(KEYINPUT96), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT97), .B(G2078), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n712), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n783), .A2(new_n771), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n784), .A2(new_n789), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n712), .A2(G4), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n632), .B2(new_n712), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1348), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n769), .A2(G26), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT28), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n466), .A2(G116), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n495), .A2(G128), .A3(new_n465), .A4(G2105), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n495), .A2(G140), .A3(new_n465), .A4(new_n466), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n802), .B1(new_n810), .B2(new_n749), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT91), .B(G2067), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G2084), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT24), .B(G34), .Z(new_n815));
  OAI22_X1  g390(.A1(new_n486), .A2(new_n749), .B1(new_n735), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n813), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n712), .A2(G21), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G168), .B2(new_n712), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G1966), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n817), .B(new_n820), .C1(new_n814), .C2(new_n816), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n712), .A2(G5), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G171), .B2(new_n712), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT95), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1961), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n797), .A2(new_n800), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n735), .A2(G35), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G162), .B2(new_n735), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT29), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2090), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n819), .A2(G1966), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT94), .Z(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n743), .A2(new_n826), .A3(new_n833), .ZN(G150));
  INV_X1    g409(.A(G150), .ZN(G311));
  NOR2_X1   g410(.A1(new_n631), .A2(new_n640), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n567), .A2(new_n571), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n534), .A2(new_n840), .B1(new_n841), .B2(new_n529), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n533), .A2(G67), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n568), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n839), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n838), .A2(new_n847), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT100), .B(G860), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n846), .A2(new_n851), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  AOI21_X1  g430(.A(new_n486), .B1(new_n499), .B2(new_n504), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n499), .A2(new_n486), .A3(new_n504), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n768), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n861));
  INV_X1    g436(.A(new_n507), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n510), .A2(new_n864), .A3(new_n515), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n510), .B2(new_n515), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n809), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n810), .B(new_n863), .C1(new_n866), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n778), .A2(new_n763), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n782), .B2(new_n764), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n495), .A2(G130), .A3(new_n465), .A4(G2105), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n495), .A2(G142), .A3(new_n465), .A4(new_n466), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT103), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n878), .A2(new_n466), .A3(G118), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(KEYINPUT103), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n466), .B2(G118), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n877), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n874), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n653), .A3(new_n652), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n654), .A2(new_n874), .A3(new_n875), .A4(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(new_n734), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n884), .A2(new_n885), .B1(new_n731), .B2(new_n733), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n763), .B1(new_n779), .B2(new_n781), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n868), .B(new_n869), .C1(new_n890), .C2(new_n871), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n873), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n860), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n873), .A2(new_n891), .ZN(new_n895));
  INV_X1    g470(.A(new_n889), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n873), .A2(new_n889), .A3(new_n891), .A4(KEYINPUT104), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n897), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(new_n903), .A3(new_n860), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n902), .B2(new_n860), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT106), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n898), .B(new_n908), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g486(.A1(new_n631), .A2(G559), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n572), .B(new_n846), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n628), .A2(new_n630), .A3(G299), .ZN(new_n915));
  AOI21_X1  g490(.A(G299), .B1(new_n628), .B2(new_n630), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n915), .B2(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n631), .A2(new_n636), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n628), .A2(new_n630), .A3(G299), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n918), .B1(new_n914), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G166), .B(G305), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n613), .B(G288), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT42), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n925), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G868), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(G868), .B2(new_n846), .ZN(G295));
  OAI21_X1  g507(.A(new_n931), .B1(G868), .B2(new_n846), .ZN(G331));
  NAND2_X1  g508(.A1(G301), .A2(KEYINPUT108), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n935), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n936));
  AND4_X1   g511(.A1(new_n553), .A2(new_n552), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n553), .A2(new_n552), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n847), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(G168), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n552), .A2(new_n934), .A3(new_n553), .A4(new_n936), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n913), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(KEYINPUT110), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n847), .B(new_n945), .C1(new_n937), .C2(new_n938), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n917), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n847), .B(new_n950), .C1(new_n937), .C2(new_n938), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n939), .A2(KEYINPUT109), .A3(new_n943), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n924), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n928), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT111), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n949), .A2(new_n953), .A3(new_n957), .A4(new_n928), .ZN(new_n958));
  INV_X1    g533(.A(new_n928), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n924), .A2(new_n951), .A3(new_n952), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n917), .B1(new_n944), .B2(new_n946), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n954), .B2(KEYINPUT111), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n947), .B1(new_n920), .B2(new_n923), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n917), .B1(new_n952), .B2(new_n951), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n959), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n965), .A2(new_n966), .A3(new_n958), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n965), .A2(new_n958), .A3(new_n969), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n973), .B1(new_n978), .B2(new_n979), .ZN(G397));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n867), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n473), .A2(G40), .A3(new_n474), .A4(new_n485), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT125), .Z(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT48), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n809), .B(G2067), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT113), .ZN(new_n991));
  INV_X1    g566(.A(new_n986), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n986), .A2(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n782), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n778), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n993), .B(new_n995), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n734), .B(new_n737), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n734), .A2(new_n737), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n998), .A2(new_n1002), .B1(G2067), .B2(new_n809), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n989), .A2(new_n1000), .B1(new_n992), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n993), .A2(KEYINPUT123), .A3(new_n997), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT123), .B1(new_n993), .B2(new_n997), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n994), .B(KEYINPUT46), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n981), .B1(new_n509), .B2(new_n516), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n984), .B1(new_n983), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G1971), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n867), .B2(new_n981), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1017), .B(new_n981), .C1(new_n509), .C2(new_n516), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n985), .A2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1018), .A2(new_n1020), .A3(G2090), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1023));
  NOR2_X1   g598(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G303), .A2(G8), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(G166), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n601), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n596), .A2(new_n597), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G651), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n599), .A2(KEYINPUT115), .A3(new_n600), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G1981), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n598), .A2(new_n601), .A3(G1981), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1032), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT116), .B1(new_n1038), .B2(G1981), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1031), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1043), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1040), .B1(new_n1038), .B2(G1981), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1045), .B(KEYINPUT49), .C1(new_n1032), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n516), .A2(KEYINPUT101), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n510), .A2(new_n515), .A3(new_n864), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n509), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G1384), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1027), .B1(new_n1051), .B2(new_n985), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1044), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT117), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1044), .A2(new_n1047), .A3(new_n1055), .A4(new_n1052), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1052), .B1(new_n1058), .B2(G288), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1052), .B(new_n1061), .C1(new_n1058), .C2(G288), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1029), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n984), .B1(KEYINPUT50), .B2(new_n1012), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n867), .A2(new_n1017), .A3(new_n981), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(G2090), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1064), .B(G8), .C1(new_n1016), .C2(new_n1068), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n1030), .A2(new_n1057), .A3(new_n1063), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1013), .A2(new_n1072), .A3(new_n1014), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1067), .A2(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1012), .A2(new_n983), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n982), .A2(new_n983), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1074), .A2(G2078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n985), .A3(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1075), .B(new_n1077), .C1(new_n1079), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1080), .A2(new_n1014), .A3(new_n985), .A4(new_n1081), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1075), .A2(new_n1077), .A3(new_n1085), .A4(G301), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1071), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1075), .A2(new_n1077), .A3(new_n1085), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1071), .B1(new_n1092), .B2(G171), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G171), .B2(new_n1083), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1080), .A2(new_n985), .A3(new_n1078), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n814), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1095), .B(G8), .C1(new_n1101), .C2(G286), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G168), .A2(new_n1027), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1097), .A2(new_n1096), .B1(new_n1099), .B2(new_n814), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1104), .B(KEYINPUT51), .C1(new_n1105), .C2(new_n1027), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1070), .A2(new_n1091), .A3(new_n1094), .A4(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1013), .A2(new_n1014), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT118), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(new_n1112), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(G299), .B(KEYINPUT57), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1118), .B(new_n1111), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT121), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT61), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n982), .A2(G2067), .A3(new_n984), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(new_n1125), .C1(new_n1099), .C2(G1348), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n982), .A2(G2067), .A3(new_n984), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n631), .B1(new_n1130), .B2(KEYINPUT60), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1132), .B(new_n632), .C1(new_n1126), .C2(new_n1129), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1131), .A2(new_n1133), .B1(KEYINPUT60), .B2(new_n1130), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT121), .B(new_n1135), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1015), .A2(new_n996), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n982), .B2(new_n984), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n839), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT59), .Z(new_n1141));
  NAND4_X1  g716(.A1(new_n1123), .A2(new_n1134), .A3(new_n1136), .A4(new_n1141), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1130), .A2(new_n631), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1121), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1143), .A2(KEYINPUT120), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT120), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1109), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1070), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1108), .A2(KEYINPUT62), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1102), .A2(new_n1106), .A3(new_n1151), .A4(new_n1107), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1084), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1105), .A2(new_n1027), .A3(G286), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1149), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1057), .A2(new_n1063), .A3(new_n1069), .ZN(new_n1159));
  OAI21_X1  g734(.A(G8), .B1(new_n1016), .B2(new_n1068), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1029), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1155), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT63), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g738(.A(G1976), .B(G288), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1052), .B1(new_n1164), .B2(new_n1040), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1163), .B(new_n1165), .C1(new_n1069), .C2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1148), .A2(new_n1158), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n613), .B(G1986), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1000), .B1(new_n986), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1011), .B1(new_n1168), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n1173));
  OR2_X1    g747(.A1(new_n460), .A2(G227), .ZN(new_n1174));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1175));
  AOI21_X1  g749(.A(G401), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g750(.A(new_n707), .B(new_n1176), .C1(new_n1175), .C2(new_n1174), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1177), .B1(new_n907), .B2(new_n909), .ZN(new_n1178));
  AND3_X1   g752(.A1(new_n971), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n1173), .B1(new_n971), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1179), .A2(new_n1180), .ZN(G308));
  NAND2_X1  g755(.A1(new_n971), .A2(new_n1178), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1182), .A2(KEYINPUT127), .ZN(new_n1183));
  NAND3_X1  g757(.A1(new_n971), .A2(new_n1178), .A3(new_n1173), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1184), .ZN(G225));
endmodule


