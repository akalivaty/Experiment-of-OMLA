

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804;

  INV_X1 U371 ( .A(n793), .ZN(n350) );
  INV_X1 U372 ( .A(G146), .ZN(n535) );
  BUF_X4 U373 ( .A(G953), .Z(n793) );
  XNOR2_X1 U374 ( .A(G116), .B(G113), .ZN(n493) );
  NOR2_X1 U375 ( .A1(n778), .A2(n666), .ZN(n769) );
  BUF_X1 U376 ( .A(n663), .Z(n778) );
  NAND2_X4 U377 ( .A1(n671), .A2(n793), .ZN(n701) );
  XNOR2_X2 U378 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X2 U379 ( .A(n690), .B(n689), .ZN(n691) );
  INV_X2 U380 ( .A(n348), .ZN(n777) );
  NAND2_X2 U381 ( .A1(n774), .A2(n349), .ZN(n348) );
  AND2_X2 U382 ( .A1(n775), .A2(n350), .ZN(n349) );
  OR2_X2 U383 ( .A1(n770), .A2(KEYINPUT2), .ZN(n771) );
  NAND2_X2 U384 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X2 U385 ( .A(n524), .B(n525), .ZN(n700) );
  XNOR2_X2 U386 ( .A(n651), .B(n650), .ZN(n655) );
  XNOR2_X2 U387 ( .A(n598), .B(n373), .ZN(n451) );
  OR2_X2 U388 ( .A1(n675), .A2(G902), .ZN(n550) );
  XNOR2_X2 U389 ( .A(n550), .B(G472), .ZN(n741) );
  NOR2_X1 U390 ( .A1(n424), .A2(KEYINPUT34), .ZN(n351) );
  AND2_X2 U391 ( .A1(n375), .A2(n376), .ZN(n367) );
  AND2_X2 U392 ( .A1(n703), .A2(G217), .ZN(n699) );
  NOR2_X2 U393 ( .A1(n449), .A2(n611), .ZN(n612) );
  INV_X1 U394 ( .A(n793), .ZN(n573) );
  XNOR2_X1 U395 ( .A(n549), .B(n541), .ZN(n410) );
  XNOR2_X1 U396 ( .A(n641), .B(KEYINPUT42), .ZN(n803) );
  XNOR2_X1 U397 ( .A(n626), .B(KEYINPUT1), .ZN(n734) );
  XNOR2_X1 U398 ( .A(n448), .B(KEYINPUT6), .ZN(n611) );
  XNOR2_X1 U399 ( .A(n549), .B(n548), .ZN(n675) );
  INV_X1 U400 ( .A(KEYINPUT45), .ZN(n467) );
  AND2_X1 U401 ( .A1(n461), .A2(n462), .ZN(n366) );
  AND2_X1 U402 ( .A1(n802), .A2(n619), .ZN(n390) );
  AND2_X1 U403 ( .A1(n398), .A2(n387), .ZN(n396) );
  AND2_X1 U404 ( .A1(n455), .A2(n454), .ZN(n453) );
  NOR2_X1 U405 ( .A1(n360), .A2(n359), .ZN(n386) );
  OR2_X1 U406 ( .A1(n451), .A2(n370), .ZN(n455) );
  NOR2_X1 U407 ( .A1(n803), .A2(KEYINPUT46), .ZN(n353) );
  NAND2_X1 U408 ( .A1(n803), .A2(KEYINPUT46), .ZN(n361) );
  XNOR2_X1 U409 ( .A(n434), .B(KEYINPUT74), .ZN(n720) );
  NOR2_X1 U410 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U411 ( .A1(n640), .A2(n629), .ZN(n434) );
  BUF_X1 U412 ( .A(n756), .Z(n766) );
  AND2_X1 U413 ( .A1(n378), .A2(n648), .ZN(n374) );
  AND2_X1 U414 ( .A1(n356), .A2(n355), .ZN(n441) );
  XNOR2_X1 U415 ( .A(n446), .B(KEYINPUT84), .ZN(n648) );
  NOR2_X1 U416 ( .A1(n610), .A2(n599), .ZN(n743) );
  XNOR2_X1 U417 ( .A(n610), .B(KEYINPUT102), .ZN(n449) );
  NAND2_X1 U418 ( .A1(n418), .A2(n413), .ZN(n368) );
  AND2_X1 U419 ( .A1(n611), .A2(n379), .ZN(n378) );
  XNOR2_X1 U420 ( .A(n502), .B(KEYINPUT38), .ZN(n749) );
  XNOR2_X1 U421 ( .A(n543), .B(n542), .ZN(n600) );
  NAND2_X1 U422 ( .A1(n734), .A2(n735), .ZN(n610) );
  BUF_X2 U423 ( .A(n734), .Z(n446) );
  AND2_X1 U424 ( .A1(n589), .A2(n603), .ZN(n747) );
  AND2_X1 U425 ( .A1(n442), .A2(n475), .ZN(n379) );
  BUF_X1 U426 ( .A(n741), .Z(n448) );
  XNOR2_X1 U427 ( .A(n741), .B(n551), .ZN(n624) );
  XNOR2_X1 U428 ( .A(n423), .B(n422), .ZN(n589) );
  AND2_X1 U429 ( .A1(n410), .A2(G469), .ZN(n362) );
  XOR2_X1 U430 ( .A(KEYINPUT62), .B(n675), .Z(n676) );
  INV_X1 U431 ( .A(n587), .ZN(n355) );
  OR2_X1 U432 ( .A1(n690), .A2(G902), .ZN(n423) );
  XNOR2_X1 U433 ( .A(n410), .B(n668), .ZN(n669) );
  XNOR2_X1 U434 ( .A(n420), .B(n365), .ZN(n570) );
  XNOR2_X1 U435 ( .A(n789), .B(n388), .ZN(n365) );
  NOR2_X1 U436 ( .A1(n793), .A2(G237), .ZN(n564) );
  XNOR2_X1 U437 ( .A(n445), .B(G104), .ZN(n538) );
  XOR2_X1 U438 ( .A(G101), .B(G140), .Z(n537) );
  XNOR2_X2 U439 ( .A(G101), .B(KEYINPUT86), .ZN(n492) );
  AND2_X1 U440 ( .A1(G902), .A2(G469), .ZN(n409) );
  XNOR2_X1 U441 ( .A(G134), .B(G116), .ZN(n554) );
  INV_X1 U442 ( .A(KEYINPUT31), .ZN(n373) );
  NAND2_X2 U443 ( .A1(n396), .A2(n394), .ZN(n802) );
  XNOR2_X1 U444 ( .A(n491), .B(n534), .ZN(n498) );
  NAND2_X1 U445 ( .A1(n386), .A2(n382), .ZN(n651) );
  XNOR2_X2 U446 ( .A(n790), .B(n535), .ZN(n549) );
  NAND2_X1 U447 ( .A1(n352), .A2(n361), .ZN(n360) );
  NAND2_X1 U448 ( .A1(n354), .A2(n353), .ZN(n352) );
  INV_X1 U449 ( .A(n801), .ZN(n354) );
  XNOR2_X2 U450 ( .A(n635), .B(n636), .ZN(n801) );
  NAND2_X1 U451 ( .A1(n358), .A2(n441), .ZN(n634) );
  XNOR2_X1 U452 ( .A(n600), .B(n357), .ZN(n356) );
  INV_X1 U453 ( .A(KEYINPUT105), .ZN(n357) );
  AND2_X2 U454 ( .A1(n458), .A2(n749), .ZN(n358) );
  XNOR2_X2 U455 ( .A(n459), .B(n473), .ZN(n458) );
  AND2_X1 U456 ( .A1(n801), .A2(KEYINPUT46), .ZN(n359) );
  NOR2_X1 U457 ( .A1(n362), .A2(n409), .ZN(n408) );
  NAND2_X1 U458 ( .A1(n377), .A2(KEYINPUT32), .ZN(n376) );
  NAND2_X1 U459 ( .A1(n466), .A2(n366), .ZN(n444) );
  XNOR2_X1 U460 ( .A(n444), .B(n467), .ZN(n663) );
  NAND2_X1 U461 ( .A1(n363), .A2(n401), .ZN(n400) );
  NAND2_X1 U462 ( .A1(n364), .A2(n351), .ZN(n363) );
  INV_X1 U463 ( .A(n756), .ZN(n364) );
  NAND2_X1 U464 ( .A1(n696), .A2(n617), .ZN(n618) );
  XNOR2_X1 U465 ( .A(n643), .B(KEYINPUT19), .ZN(n628) );
  NAND2_X1 U466 ( .A1(n380), .A2(n367), .ZN(n696) );
  NOR2_X1 U467 ( .A1(n628), .A2(n385), .ZN(n440) );
  NAND2_X2 U468 ( .A1(n369), .A2(n368), .ZN(n643) );
  AND2_X2 U469 ( .A1(n415), .A2(n414), .ZN(n369) );
  INV_X1 U470 ( .A(KEYINPUT95), .ZN(n370) );
  OR2_X1 U471 ( .A1(n451), .A2(n371), .ZN(n724) );
  INV_X1 U472 ( .A(n723), .ZN(n371) );
  OR2_X1 U473 ( .A1(n451), .A2(n372), .ZN(n726) );
  INV_X1 U474 ( .A(n725), .ZN(n372) );
  NAND2_X1 U475 ( .A1(n605), .A2(n374), .ZN(n375) );
  NAND2_X1 U476 ( .A1(n648), .A2(n442), .ZN(n377) );
  NAND2_X1 U477 ( .A1(n605), .A2(n611), .ZN(n616) );
  NAND2_X1 U478 ( .A1(n616), .A2(KEYINPUT32), .ZN(n380) );
  XNOR2_X2 U479 ( .A(n618), .B(n438), .ZN(n435) );
  NAND2_X1 U480 ( .A1(n482), .A2(n476), .ZN(n381) );
  NAND2_X1 U481 ( .A1(n482), .A2(n476), .ZN(n417) );
  XNOR2_X2 U482 ( .A(n580), .B(KEYINPUT22), .ZN(n605) );
  XNOR2_X2 U483 ( .A(n498), .B(n783), .ZN(n681) );
  INV_X1 U484 ( .A(n613), .ZN(n597) );
  XNOR2_X1 U485 ( .A(n571), .B(G475), .ZN(n422) );
  XNOR2_X1 U486 ( .A(KEYINPUT10), .B(G140), .ZN(n518) );
  INV_X1 U487 ( .A(KEYINPUT99), .ZN(n456) );
  XNOR2_X1 U488 ( .A(G902), .B(KEYINPUT15), .ZN(n507) );
  NOR2_X1 U489 ( .A1(n477), .A2(n483), .ZN(n476) );
  XNOR2_X1 U490 ( .A(G131), .B(G134), .ZN(n531) );
  XOR2_X1 U491 ( .A(G137), .B(KEYINPUT67), .Z(n532) );
  AND2_X1 U492 ( .A1(n402), .A2(n614), .ZN(n401) );
  NOR2_X1 U493 ( .A1(n577), .A2(n506), .ZN(n587) );
  NAND2_X2 U494 ( .A1(n408), .A2(n404), .ZN(n626) );
  NAND2_X1 U495 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U496 ( .A(n530), .B(n529), .ZN(n731) );
  XNOR2_X1 U497 ( .A(KEYINPUT16), .B(G122), .ZN(n496) );
  XNOR2_X1 U498 ( .A(n522), .B(n443), .ZN(n553) );
  XNOR2_X1 U499 ( .A(n523), .B(n521), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n570), .B(n569), .ZN(n690) );
  XNOR2_X1 U501 ( .A(G143), .B(G131), .ZN(n567) );
  NOR2_X1 U502 ( .A1(n397), .A2(n403), .ZN(n393) );
  INV_X1 U503 ( .A(n400), .ZN(n395) );
  INV_X1 U504 ( .A(KEYINPUT30), .ZN(n473) );
  INV_X1 U505 ( .A(KEYINPUT82), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n435), .B(n437), .ZN(n436) );
  INV_X1 U507 ( .A(KEYINPUT81), .ZN(n437) );
  INV_X1 U508 ( .A(n728), .ZN(n447) );
  INV_X1 U509 ( .A(KEYINPUT100), .ZN(n463) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n609) );
  INV_X1 U511 ( .A(G237), .ZN(n499) );
  NAND2_X1 U512 ( .A1(n501), .A2(n658), .ZN(n481) );
  NAND2_X1 U513 ( .A1(n480), .A2(n507), .ZN(n479) );
  INV_X1 U514 ( .A(n501), .ZN(n480) );
  NAND2_X1 U515 ( .A1(n416), .A2(KEYINPUT83), .ZN(n414) );
  INV_X1 U516 ( .A(n478), .ZN(n416) );
  INV_X1 U517 ( .A(G469), .ZN(n407) );
  XNOR2_X1 U518 ( .A(KEYINPUT3), .B(G119), .ZN(n494) );
  XNOR2_X1 U519 ( .A(n421), .B(KEYINPUT97), .ZN(n420) );
  NAND2_X1 U520 ( .A1(n564), .A2(G214), .ZN(n421) );
  XNOR2_X1 U521 ( .A(G113), .B(G104), .ZN(n565) );
  XOR2_X1 U522 ( .A(KEYINPUT11), .B(G122), .Z(n566) );
  NAND2_X1 U523 ( .A1(G234), .A2(G237), .ZN(n503) );
  XNOR2_X1 U524 ( .A(n440), .B(n439), .ZN(n613) );
  INV_X1 U525 ( .A(KEYINPUT0), .ZN(n439) );
  BUF_X1 U526 ( .A(n664), .Z(n796) );
  XOR2_X1 U527 ( .A(G122), .B(G107), .Z(n555) );
  INV_X1 U528 ( .A(KEYINPUT32), .ZN(n475) );
  XNOR2_X1 U529 ( .A(n465), .B(n464), .ZN(n627) );
  INV_X1 U530 ( .A(KEYINPUT28), .ZN(n464) );
  INV_X1 U531 ( .A(KEYINPUT94), .ZN(n542) );
  BUF_X1 U532 ( .A(n731), .Z(n442) );
  XNOR2_X1 U533 ( .A(n520), .B(n789), .ZN(n525) );
  NAND2_X1 U534 ( .A1(n427), .A2(n428), .ZN(n430) );
  INV_X1 U535 ( .A(KEYINPUT78), .ZN(n428) );
  NAND2_X1 U536 ( .A1(n395), .A2(n392), .ZN(n394) );
  INV_X1 U537 ( .A(n614), .ZN(n411) );
  NOR2_X1 U538 ( .A1(n642), .A2(n447), .ZN(n382) );
  AND2_X1 U539 ( .A1(n713), .A2(KEYINPUT95), .ZN(n383) );
  AND2_X1 U540 ( .A1(n802), .A2(KEYINPUT69), .ZN(n384) );
  XNOR2_X1 U541 ( .A(n578), .B(KEYINPUT90), .ZN(n385) );
  NAND2_X1 U542 ( .A1(n766), .A2(n393), .ZN(n387) );
  XNOR2_X1 U543 ( .A(KEYINPUT12), .B(KEYINPUT96), .ZN(n388) );
  AND2_X1 U544 ( .A1(n802), .A2(n474), .ZN(n389) );
  INV_X1 U545 ( .A(KEYINPUT83), .ZN(n419) );
  AND2_X1 U546 ( .A1(n478), .A2(n481), .ZN(n391) );
  AND2_X1 U547 ( .A1(n399), .A2(n397), .ZN(n392) );
  INV_X1 U548 ( .A(G902), .ZN(n406) );
  NAND2_X1 U549 ( .A1(n756), .A2(KEYINPUT34), .ZN(n399) );
  INV_X1 U550 ( .A(n615), .ZN(n397) );
  NAND2_X1 U551 ( .A1(n400), .A2(n615), .ZN(n398) );
  NAND2_X1 U552 ( .A1(n424), .A2(KEYINPUT34), .ZN(n402) );
  INV_X1 U553 ( .A(KEYINPUT34), .ZN(n403) );
  OR2_X1 U554 ( .A1(n410), .A2(n405), .ZN(n404) );
  NAND2_X1 U555 ( .A1(n441), .A2(n458), .ZN(n412) );
  NOR2_X1 U556 ( .A1(n412), .A2(n411), .ZN(n572) );
  INV_X1 U557 ( .A(n381), .ZN(n413) );
  NAND2_X1 U558 ( .A1(n417), .A2(KEYINPUT83), .ZN(n415) );
  AND2_X1 U559 ( .A1(n478), .A2(n419), .ZN(n418) );
  INV_X1 U560 ( .A(n597), .ZN(n424) );
  NAND2_X1 U561 ( .A1(n391), .A2(n482), .ZN(n502) );
  BUF_X1 U562 ( .A(n559), .Z(n425) );
  BUF_X1 U563 ( .A(n790), .Z(n426) );
  NAND2_X1 U564 ( .A1(n773), .A2(KEYINPUT78), .ZN(n429) );
  NAND2_X1 U565 ( .A1(n429), .A2(n430), .ZN(n774) );
  INV_X1 U566 ( .A(n773), .ZN(n427) );
  BUF_X1 U567 ( .A(n801), .Z(n431) );
  NAND2_X1 U568 ( .A1(n432), .A2(n633), .ZN(n642) );
  NAND2_X1 U569 ( .A1(n632), .A2(n631), .ZN(n432) );
  XNOR2_X1 U570 ( .A(n433), .B(KEYINPUT103), .ZN(n590) );
  NAND2_X1 U571 ( .A1(n588), .A2(n625), .ZN(n433) );
  NAND2_X1 U572 ( .A1(n390), .A2(n435), .ZN(n460) );
  NAND2_X1 U573 ( .A1(n436), .A2(n389), .ZN(n471) );
  NAND2_X1 U574 ( .A1(n436), .A2(n384), .ZN(n469) );
  XNOR2_X1 U575 ( .A(n634), .B(KEYINPUT39), .ZN(n652) );
  XNOR2_X2 U576 ( .A(G110), .B(G107), .ZN(n445) );
  NAND2_X1 U577 ( .A1(n626), .A2(n735), .ZN(n543) );
  NAND2_X1 U578 ( .A1(n652), .A2(n723), .ZN(n635) );
  NAND2_X1 U579 ( .A1(n470), .A2(n469), .ZN(n466) );
  NAND2_X1 U580 ( .A1(n451), .A2(n450), .ZN(n454) );
  NOR2_X1 U581 ( .A1(n713), .A2(KEYINPUT95), .ZN(n450) );
  NAND2_X1 U582 ( .A1(n453), .A2(n452), .ZN(n457) );
  NOR2_X1 U583 ( .A1(n383), .A2(n630), .ZN(n452) );
  XNOR2_X2 U584 ( .A(n534), .B(n533), .ZN(n790) );
  NAND2_X1 U585 ( .A1(n624), .A2(n748), .ZN(n459) );
  XNOR2_X1 U586 ( .A(n468), .B(n463), .ZN(n461) );
  NAND2_X1 U587 ( .A1(n460), .A2(KEYINPUT44), .ZN(n462) );
  NAND2_X1 U588 ( .A1(n624), .A2(n625), .ZN(n465) );
  NAND2_X1 U589 ( .A1(n609), .A2(n710), .ZN(n468) );
  NAND2_X1 U590 ( .A1(n471), .A2(n619), .ZN(n470) );
  NAND2_X1 U591 ( .A1(n597), .A2(n743), .ZN(n598) );
  XNOR2_X2 U592 ( .A(n472), .B(G143), .ZN(n559) );
  XNOR2_X2 U593 ( .A(G128), .B(KEYINPUT64), .ZN(n472) );
  INV_X1 U594 ( .A(KEYINPUT44), .ZN(n474) );
  INV_X1 U595 ( .A(n481), .ZN(n477) );
  OR2_X2 U596 ( .A1(n681), .A2(n479), .ZN(n478) );
  NAND2_X1 U597 ( .A1(n681), .A2(n501), .ZN(n482) );
  INV_X1 U598 ( .A(n748), .ZN(n483) );
  BUF_X1 U599 ( .A(n698), .Z(n703) );
  INV_X1 U600 ( .A(n630), .ZN(n604) );
  INV_X1 U601 ( .A(KEYINPUT77), .ZN(n521) );
  INV_X1 U602 ( .A(G953), .ZN(n484) );
  NAND2_X1 U603 ( .A1(n484), .A2(G224), .ZN(n485) );
  XNOR2_X1 U604 ( .A(n485), .B(KEYINPUT72), .ZN(n486) );
  XNOR2_X1 U605 ( .A(G146), .B(G125), .ZN(n519) );
  XNOR2_X1 U606 ( .A(n486), .B(n519), .ZN(n490) );
  XNOR2_X1 U607 ( .A(KEYINPUT87), .B(KEYINPUT17), .ZN(n488) );
  XNOR2_X1 U608 ( .A(KEYINPUT18), .B(KEYINPUT73), .ZN(n487) );
  XNOR2_X1 U609 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U610 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X2 U611 ( .A(n559), .B(KEYINPUT4), .ZN(n534) );
  XNOR2_X1 U612 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X2 U613 ( .A(n495), .B(n494), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n538), .B(n496), .ZN(n497) );
  XNOR2_X2 U615 ( .A(n547), .B(n497), .ZN(n783) );
  INV_X1 U616 ( .A(n507), .ZN(n658) );
  NAND2_X1 U617 ( .A1(n406), .A2(n499), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n552), .A2(G210), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n500), .B(KEYINPUT88), .ZN(n501) );
  INV_X1 U620 ( .A(n502), .ZN(n595) );
  XNOR2_X1 U621 ( .A(n503), .B(KEYINPUT14), .ZN(n504) );
  NAND2_X1 U622 ( .A1(G952), .A2(n504), .ZN(n763) );
  NOR2_X1 U623 ( .A1(n793), .A2(n763), .ZN(n577) );
  AND2_X1 U624 ( .A1(G902), .A2(n504), .ZN(n574) );
  NAND2_X1 U625 ( .A1(n793), .A2(n574), .ZN(n505) );
  NOR2_X1 U626 ( .A1(G900), .A2(n505), .ZN(n506) );
  NAND2_X1 U627 ( .A1(G234), .A2(n507), .ZN(n508) );
  XNOR2_X1 U628 ( .A(KEYINPUT20), .B(n508), .ZN(n526) );
  NAND2_X1 U629 ( .A1(G221), .A2(n526), .ZN(n511) );
  INV_X1 U630 ( .A(KEYINPUT93), .ZN(n509) );
  XNOR2_X1 U631 ( .A(n509), .B(KEYINPUT21), .ZN(n510) );
  XNOR2_X1 U632 ( .A(n511), .B(n510), .ZN(n730) );
  XOR2_X1 U633 ( .A(G110), .B(G119), .Z(n513) );
  XNOR2_X1 U634 ( .A(G128), .B(G137), .ZN(n512) );
  XNOR2_X1 U635 ( .A(n513), .B(n512), .ZN(n517) );
  XOR2_X1 U636 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n515) );
  XNOR2_X1 U637 ( .A(KEYINPUT91), .B(KEYINPUT23), .ZN(n514) );
  XNOR2_X1 U638 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U639 ( .A(n517), .B(n516), .ZN(n520) );
  XNOR2_X1 U640 ( .A(n519), .B(n518), .ZN(n789) );
  AND2_X1 U641 ( .A1(G234), .A2(n573), .ZN(n522) );
  XNOR2_X1 U642 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n523) );
  NAND2_X1 U643 ( .A1(G221), .A2(n553), .ZN(n524) );
  NAND2_X1 U644 ( .A1(n700), .A2(n406), .ZN(n530) );
  NAND2_X1 U645 ( .A1(n526), .A2(G217), .ZN(n527) );
  XNOR2_X1 U646 ( .A(n527), .B(KEYINPUT71), .ZN(n528) );
  XOR2_X1 U647 ( .A(KEYINPUT25), .B(n528), .Z(n529) );
  NOR2_X2 U648 ( .A1(n730), .A2(n731), .ZN(n735) );
  XNOR2_X1 U649 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U650 ( .A1(G227), .A2(n573), .ZN(n536) );
  XNOR2_X1 U651 ( .A(n537), .B(n536), .ZN(n540) );
  INV_X1 U652 ( .A(n538), .ZN(n539) );
  XNOR2_X1 U653 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U654 ( .A(KEYINPUT70), .B(KEYINPUT5), .Z(n545) );
  NAND2_X1 U655 ( .A1(n564), .A2(G210), .ZN(n544) );
  XNOR2_X1 U656 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U657 ( .A(n547), .B(n546), .ZN(n548) );
  INV_X1 U658 ( .A(KEYINPUT101), .ZN(n551) );
  NAND2_X1 U659 ( .A1(n552), .A2(G214), .ZN(n748) );
  NAND2_X1 U660 ( .A1(G217), .A2(n553), .ZN(n557) );
  XNOR2_X1 U661 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U662 ( .A(n557), .B(n556), .ZN(n561) );
  XNOR2_X1 U663 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n558) );
  XNOR2_X1 U664 ( .A(n425), .B(n558), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n561), .B(n560), .ZN(n704) );
  NAND2_X1 U666 ( .A1(n704), .A2(n406), .ZN(n563) );
  INV_X1 U667 ( .A(G478), .ZN(n562) );
  XNOR2_X1 U668 ( .A(n563), .B(n562), .ZN(n603) );
  XNOR2_X1 U669 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n571) );
  XNOR2_X1 U670 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U671 ( .A(n568), .B(n567), .Z(n569) );
  NOR2_X1 U672 ( .A1(n603), .A2(n589), .ZN(n614) );
  NAND2_X1 U673 ( .A1(n595), .A2(n572), .ZN(n621) );
  XNOR2_X1 U674 ( .A(n621), .B(G143), .ZN(G45) );
  NOR2_X1 U675 ( .A1(G898), .A2(n573), .ZN(n784) );
  NAND2_X1 U676 ( .A1(n574), .A2(n784), .ZN(n575) );
  XNOR2_X1 U677 ( .A(KEYINPUT89), .B(n575), .ZN(n576) );
  NOR2_X1 U678 ( .A1(n577), .A2(n576), .ZN(n578) );
  INV_X1 U679 ( .A(n730), .ZN(n585) );
  NAND2_X1 U680 ( .A1(n747), .A2(n585), .ZN(n579) );
  NOR2_X2 U681 ( .A1(n613), .A2(n579), .ZN(n580) );
  BUF_X1 U682 ( .A(n605), .Z(n584) );
  INV_X1 U683 ( .A(n442), .ZN(n581) );
  OR2_X1 U684 ( .A1(n446), .A2(n581), .ZN(n582) );
  NOR2_X1 U685 ( .A1(n582), .A2(n624), .ZN(n583) );
  NAND2_X1 U686 ( .A1(n584), .A2(n583), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(G110), .ZN(G12) );
  XNOR2_X1 U688 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n594) );
  INV_X1 U689 ( .A(n611), .ZN(n588) );
  NAND2_X1 U690 ( .A1(n731), .A2(n585), .ZN(n586) );
  NOR2_X1 U691 ( .A1(n587), .A2(n586), .ZN(n625) );
  INV_X1 U692 ( .A(n589), .ZN(n602) );
  AND2_X1 U693 ( .A1(n603), .A2(n602), .ZN(n723) );
  NAND2_X1 U694 ( .A1(n590), .A2(n723), .ZN(n646) );
  INV_X1 U695 ( .A(n646), .ZN(n591) );
  NAND2_X1 U696 ( .A1(n591), .A2(n748), .ZN(n592) );
  NOR2_X1 U697 ( .A1(n446), .A2(n592), .ZN(n593) );
  XNOR2_X1 U698 ( .A(n594), .B(n593), .ZN(n596) );
  NOR2_X1 U699 ( .A1(n596), .A2(n595), .ZN(n653) );
  XOR2_X1 U700 ( .A(G140), .B(n653), .Z(G42) );
  INV_X1 U701 ( .A(KEYINPUT65), .ZN(n662) );
  INV_X1 U702 ( .A(n448), .ZN(n599) );
  NAND2_X1 U703 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U704 ( .A1(n424), .A2(n601), .ZN(n713) );
  NOR2_X1 U705 ( .A1(n603), .A2(n602), .ZN(n725) );
  NOR2_X1 U706 ( .A1(n723), .A2(n725), .ZN(n630) );
  BUF_X1 U707 ( .A(n616), .Z(n606) );
  XOR2_X1 U708 ( .A(KEYINPUT80), .B(n606), .Z(n608) );
  NOR2_X1 U709 ( .A1(n446), .A2(n442), .ZN(n607) );
  NAND2_X1 U710 ( .A1(n608), .A2(n607), .ZN(n710) );
  XNOR2_X1 U711 ( .A(n612), .B(KEYINPUT33), .ZN(n756) );
  XNOR2_X1 U712 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n615) );
  INV_X1 U713 ( .A(KEYINPUT69), .ZN(n619) );
  NAND2_X1 U714 ( .A1(KEYINPUT47), .A2(n630), .ZN(n620) );
  XNOR2_X1 U715 ( .A(n620), .B(KEYINPUT76), .ZN(n622) );
  NAND2_X1 U716 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U717 ( .A(KEYINPUT75), .B(n623), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n627), .A2(n626), .ZN(n640) );
  BUF_X1 U719 ( .A(n628), .Z(n629) );
  XOR2_X1 U720 ( .A(KEYINPUT47), .B(n720), .Z(n632) );
  OR2_X1 U721 ( .A1(KEYINPUT47), .A2(n604), .ZN(n631) );
  XOR2_X1 U722 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n636) );
  XOR2_X1 U723 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n639) );
  NAND2_X1 U724 ( .A1(n749), .A2(n748), .ZN(n637) );
  XNOR2_X1 U725 ( .A(n637), .B(KEYINPUT107), .ZN(n752) );
  NAND2_X1 U726 ( .A1(n752), .A2(n747), .ZN(n638) );
  XNOR2_X1 U727 ( .A(n639), .B(n638), .ZN(n765) );
  NOR2_X1 U728 ( .A1(n640), .A2(n765), .ZN(n641) );
  BUF_X1 U729 ( .A(n643), .Z(n644) );
  INV_X1 U730 ( .A(n644), .ZN(n645) );
  XNOR2_X1 U731 ( .A(n647), .B(KEYINPUT36), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n728) );
  XOR2_X1 U733 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n650) );
  AND2_X1 U734 ( .A1(n652), .A2(n725), .ZN(n729) );
  NOR2_X1 U735 ( .A1(n653), .A2(n729), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n664) );
  INV_X1 U737 ( .A(n664), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n656), .A2(n658), .ZN(n657) );
  NOR2_X1 U739 ( .A1(n663), .A2(n657), .ZN(n660) );
  AND2_X1 U740 ( .A1(n658), .A2(KEYINPUT2), .ZN(n659) );
  NOR2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(n662), .ZN(n667) );
  INV_X1 U743 ( .A(n796), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(KEYINPUT2), .ZN(n666) );
  NOR2_X2 U745 ( .A1(n667), .A2(n769), .ZN(n698) );
  NAND2_X1 U746 ( .A1(n698), .A2(G469), .ZN(n670) );
  XNOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n672) );
  INV_X1 U749 ( .A(G952), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n672), .A2(n701), .ZN(n674) );
  INV_X1 U751 ( .A(KEYINPUT120), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n674), .B(n673), .ZN(G54) );
  NAND2_X1 U753 ( .A1(n698), .A2(G472), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n678), .A2(n701), .ZN(n680) );
  XOR2_X1 U756 ( .A(KEYINPUT85), .B(KEYINPUT63), .Z(n679) );
  XNOR2_X1 U757 ( .A(n680), .B(n679), .ZN(G57) );
  NAND2_X1 U758 ( .A1(n698), .A2(G210), .ZN(n685) );
  BUF_X1 U759 ( .A(n681), .Z(n683) );
  XNOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n682) );
  XNOR2_X1 U761 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U762 ( .A1(n686), .A2(n701), .ZN(n688) );
  XNOR2_X1 U763 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n687) );
  XNOR2_X1 U764 ( .A(n688), .B(n687), .ZN(G51) );
  NAND2_X1 U765 ( .A1(n698), .A2(G475), .ZN(n692) );
  XOR2_X1 U766 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n689) );
  XNOR2_X1 U767 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n693), .A2(n701), .ZN(n695) );
  INV_X1 U769 ( .A(KEYINPUT60), .ZN(n694) );
  XNOR2_X1 U770 ( .A(n695), .B(n694), .ZN(G60) );
  BUF_X1 U771 ( .A(n696), .Z(n697) );
  XNOR2_X1 U772 ( .A(n697), .B(G119), .ZN(G21) );
  XNOR2_X1 U773 ( .A(n699), .B(n700), .ZN(n702) );
  INV_X1 U774 ( .A(n701), .ZN(n707) );
  NOR2_X1 U775 ( .A1(n702), .A2(n707), .ZN(G66) );
  NAND2_X1 U776 ( .A1(n703), .A2(G478), .ZN(n706) );
  XOR2_X1 U777 ( .A(KEYINPUT122), .B(n704), .Z(n705) );
  XNOR2_X1 U778 ( .A(n706), .B(n705), .ZN(n708) );
  NOR2_X1 U779 ( .A1(n708), .A2(n707), .ZN(G63) );
  XOR2_X1 U780 ( .A(G101), .B(KEYINPUT109), .Z(n709) );
  XNOR2_X1 U781 ( .A(n710), .B(n709), .ZN(G3) );
  NAND2_X1 U782 ( .A1(n713), .A2(n723), .ZN(n711) );
  XNOR2_X1 U783 ( .A(n711), .B(KEYINPUT110), .ZN(n712) );
  XNOR2_X1 U784 ( .A(G104), .B(n712), .ZN(G6) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n715) );
  NAND2_X1 U786 ( .A1(n713), .A2(n725), .ZN(n714) );
  XNOR2_X1 U787 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U788 ( .A(G107), .B(n716), .ZN(G9) );
  XOR2_X1 U789 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n718) );
  NAND2_X1 U790 ( .A1(n725), .A2(n720), .ZN(n717) );
  XNOR2_X1 U791 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U792 ( .A(G128), .B(n719), .Z(G30) );
  NAND2_X1 U793 ( .A1(n720), .A2(n723), .ZN(n721) );
  XNOR2_X1 U794 ( .A(n721), .B(KEYINPUT112), .ZN(n722) );
  XNOR2_X1 U795 ( .A(G146), .B(n722), .ZN(G48) );
  XNOR2_X1 U796 ( .A(n724), .B(G113), .ZN(G15) );
  XNOR2_X1 U797 ( .A(n726), .B(G116), .ZN(G18) );
  XOR2_X1 U798 ( .A(G125), .B(KEYINPUT37), .Z(n727) );
  XNOR2_X1 U799 ( .A(n728), .B(n727), .ZN(G27) );
  XOR2_X1 U800 ( .A(G134), .B(n729), .Z(G36) );
  NAND2_X1 U801 ( .A1(n442), .A2(n730), .ZN(n732) );
  XNOR2_X1 U802 ( .A(n732), .B(KEYINPUT49), .ZN(n733) );
  XNOR2_X1 U803 ( .A(KEYINPUT113), .B(n733), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n735), .A2(n446), .ZN(n736) );
  XOR2_X1 U805 ( .A(KEYINPUT50), .B(n736), .Z(n737) );
  XNOR2_X1 U806 ( .A(KEYINPUT114), .B(n737), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U808 ( .A1(n448), .A2(n740), .ZN(n742) );
  NOR2_X1 U809 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U810 ( .A(n744), .B(KEYINPUT115), .ZN(n745) );
  XNOR2_X1 U811 ( .A(KEYINPUT51), .B(n745), .ZN(n746) );
  NOR2_X1 U812 ( .A1(n765), .A2(n746), .ZN(n759) );
  INV_X1 U813 ( .A(n747), .ZN(n751) );
  NOR2_X1 U814 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U815 ( .A1(n751), .A2(n750), .ZN(n755) );
  NAND2_X1 U816 ( .A1(n752), .A2(n604), .ZN(n753) );
  XOR2_X1 U817 ( .A(KEYINPUT116), .B(n753), .Z(n754) );
  NOR2_X1 U818 ( .A1(n755), .A2(n754), .ZN(n757) );
  NOR2_X1 U819 ( .A1(n757), .A2(n766), .ZN(n758) );
  NOR2_X1 U820 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U821 ( .A(n760), .B(KEYINPUT52), .Z(n761) );
  XNOR2_X1 U822 ( .A(KEYINPUT117), .B(n761), .ZN(n762) );
  NOR2_X1 U823 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U824 ( .A(n764), .B(KEYINPUT118), .ZN(n768) );
  NOR2_X1 U825 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U826 ( .A1(n768), .A2(n767), .ZN(n775) );
  INV_X1 U827 ( .A(n769), .ZN(n772) );
  NOR2_X1 U828 ( .A1(n778), .A2(n796), .ZN(n770) );
  XNOR2_X1 U829 ( .A(n777), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U830 ( .A1(n778), .A2(n793), .ZN(n782) );
  NAND2_X1 U831 ( .A1(n793), .A2(G224), .ZN(n779) );
  XNOR2_X1 U832 ( .A(KEYINPUT61), .B(n779), .ZN(n780) );
  AND2_X1 U833 ( .A1(n780), .A2(G898), .ZN(n781) );
  NOR2_X1 U834 ( .A1(n782), .A2(n781), .ZN(n788) );
  XOR2_X1 U835 ( .A(KEYINPUT123), .B(n783), .Z(n785) );
  NOR2_X1 U836 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U837 ( .A(KEYINPUT124), .B(n786), .Z(n787) );
  XNOR2_X1 U838 ( .A(n788), .B(n787), .ZN(G69) );
  XNOR2_X1 U839 ( .A(n426), .B(n789), .ZN(n795) );
  XOR2_X1 U840 ( .A(G227), .B(n795), .Z(n791) );
  NAND2_X1 U841 ( .A1(n791), .A2(G900), .ZN(n792) );
  NAND2_X1 U842 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U843 ( .A(n794), .B(KEYINPUT126), .ZN(n800) );
  XNOR2_X1 U844 ( .A(KEYINPUT125), .B(n795), .ZN(n797) );
  XNOR2_X1 U845 ( .A(n797), .B(n796), .ZN(n798) );
  NAND2_X1 U846 ( .A1(n798), .A2(n573), .ZN(n799) );
  NAND2_X1 U847 ( .A1(n800), .A2(n799), .ZN(G72) );
  XOR2_X1 U848 ( .A(n431), .B(G131), .Z(G33) );
  XNOR2_X1 U849 ( .A(n802), .B(G122), .ZN(G24) );
  XNOR2_X1 U850 ( .A(G137), .B(KEYINPUT127), .ZN(n804) );
  XNOR2_X1 U851 ( .A(n804), .B(n803), .ZN(G39) );
endmodule

