//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT0), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT0), .B(G128), .Z(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n189), .B2(new_n193), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT78), .A2(G107), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT78), .A2(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(G104), .A3(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(G104), .A2(G107), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT3), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n199), .A2(new_n200), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n200), .B1(new_n199), .B2(new_n204), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NOR4_X1   g023(.A1(new_n199), .A2(new_n200), .A3(new_n204), .A4(new_n207), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n194), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(G137), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT11), .A3(G134), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n214), .A2(new_n217), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n215), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n214), .A2(new_n217), .A3(new_n222), .A4(new_n215), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n195), .A2(new_n196), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n228), .B2(new_n202), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n189), .A2(new_n231), .A3(G128), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n191), .A2(new_n233), .A3(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(G146), .C1(new_n191), .C2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(KEYINPUT10), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n206), .A2(new_n237), .A3(new_n229), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n211), .A2(new_n226), .A3(new_n238), .A4(new_n241), .ZN(new_n242));
  XOR2_X1   g056(.A(G110), .B(G140), .Z(new_n243));
  INV_X1    g057(.A(G953), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n244), .A2(G227), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n243), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n206), .A2(new_n229), .ZN(new_n248));
  INV_X1    g062(.A(new_n237), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n239), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n218), .A2(G131), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT12), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n257), .B(new_n226), .C1(new_n250), .C2(new_n239), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n206), .A2(new_n208), .ZN(new_n261));
  INV_X1    g075(.A(new_n205), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n210), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n194), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n238), .B(new_n241), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n246), .B1(new_n266), .B2(new_n242), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n187), .B(new_n188), .C1(new_n260), .C2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n242), .A3(new_n246), .ZN(new_n269));
  INV_X1    g083(.A(new_n242), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(G469), .B(new_n269), .C1(new_n271), .C2(new_n246), .ZN(new_n272));
  NAND2_X1  g086(.A1(G469), .A2(G902), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G221), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT9), .B(G234), .Z(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n188), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G475), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT71), .A2(G125), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(G140), .ZN(new_n283));
  INV_X1    g097(.A(G140), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT72), .B1(new_n284), .B2(G125), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT71), .A3(G125), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n287), .A2(KEYINPUT16), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT16), .B1(new_n284), .B2(G125), .ZN(new_n289));
  OAI21_X1  g103(.A(G146), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n287), .B2(KEYINPUT16), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(new_n233), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n291), .B(G146), .C1(new_n288), .C2(new_n289), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G237), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n244), .A3(G214), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n235), .ZN(new_n300));
  NOR2_X1   g114(.A1(G237), .A2(G953), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(G214), .C1(KEYINPUT84), .C2(G143), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G131), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT17), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(new_n222), .A3(new_n302), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT88), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n304), .A2(KEYINPUT88), .A3(new_n305), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(KEYINPUT17), .A3(G131), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT87), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n296), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(new_n201), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n287), .A2(G146), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n284), .A2(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n284), .A2(G125), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n233), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(new_n322), .B(KEYINPUT85), .Z(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n303), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n315), .A2(new_n317), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n287), .A2(KEYINPUT19), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT19), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n329), .A3(new_n320), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n233), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n290), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n304), .A2(new_n306), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n290), .A2(KEYINPUT86), .A3(new_n331), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n317), .B1(new_n337), .B2(new_n326), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n280), .B(new_n188), .C1(new_n327), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n315), .A2(new_n317), .A3(new_n326), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n337), .A2(new_n326), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n317), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n344), .A2(KEYINPUT20), .A3(new_n280), .A4(new_n188), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n317), .B1(new_n315), .B2(new_n326), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n188), .B1(new_n327), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G475), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n341), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT89), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n341), .A2(new_n345), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G478), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  XNOR2_X1  g169(.A(G116), .B(G122), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n227), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT90), .ZN(new_n358));
  XNOR2_X1  g172(.A(G128), .B(G143), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(new_n213), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT14), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT14), .A3(G122), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(G107), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n213), .ZN(new_n367));
  INV_X1    g181(.A(new_n357), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n227), .A2(new_n356), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n191), .A2(KEYINPUT13), .A3(G143), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n213), .B(new_n371), .C1(KEYINPUT13), .C2(new_n359), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n358), .A2(new_n366), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n276), .A2(G217), .A3(new_n244), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n188), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT91), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n355), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n380), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(KEYINPUT91), .A3(new_n188), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n384), .B2(new_n355), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n244), .A2(G952), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(G234), .B2(G237), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT21), .B(G898), .Z(new_n389));
  NAND2_X1  g203(.A1(G234), .A2(G237), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(G902), .A3(G953), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AND4_X1   g206(.A1(new_n279), .A2(new_n353), .A3(new_n385), .A4(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n215), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n213), .A2(G137), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(new_n237), .C1(new_n253), .C2(new_n254), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(KEYINPUT30), .C1(new_n226), .C2(new_n264), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT67), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n255), .A2(new_n194), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT67), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT30), .A4(new_n397), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT65), .B1(new_n226), .B2(new_n264), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n255), .A2(new_n405), .A3(new_n194), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n397), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G116), .B(G119), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT2), .B(G113), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT2), .B(G113), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n410), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT66), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT66), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n403), .A2(new_n409), .A3(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT26), .B(G101), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n301), .A2(G210), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n400), .A2(new_n418), .A3(new_n397), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT31), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n407), .A2(new_n419), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n429), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n425), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT31), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n420), .A2(new_n436), .A3(new_n425), .A4(new_n426), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G472), .A2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT32), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n442), .A3(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n433), .A2(KEYINPUT29), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT29), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT69), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n432), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n400), .A2(new_n397), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n419), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n429), .B1(new_n450), .B2(new_n426), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT69), .B1(new_n426), .B2(new_n429), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n445), .B(new_n425), .C1(new_n446), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n420), .A2(new_n426), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n425), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n454), .B(new_n188), .C1(KEYINPUT29), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G472), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(G234), .B2(new_n188), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G119), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n463), .A2(KEYINPUT23), .A3(G128), .ZN(new_n464));
  XNOR2_X1  g278(.A(G119), .B(G128), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(KEYINPUT23), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT70), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n191), .B2(G119), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(KEYINPUT70), .A3(G128), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n468), .A2(new_n469), .B1(G119), .B2(new_n191), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT24), .B(G110), .Z(new_n471));
  AOI22_X1  g285(.A1(new_n466), .A2(G110), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n294), .A2(new_n472), .A3(new_n295), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT74), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n321), .B1(new_n292), .B2(new_n233), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT75), .B(G110), .Z(new_n477));
  OAI22_X1  g291(.A1(new_n466), .A2(new_n477), .B1(new_n470), .B2(new_n471), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n475), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n290), .A2(KEYINPUT76), .A3(new_n478), .A4(new_n321), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n294), .A2(new_n483), .A3(new_n472), .A4(new_n295), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n244), .A2(G221), .A3(G234), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT22), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(G137), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n474), .A2(new_n482), .A3(new_n484), .A4(new_n488), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n188), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n490), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n491), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n462), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n492), .A2(new_n461), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT77), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n461), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT77), .ZN(new_n501));
  INV_X1    g315(.A(new_n497), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n444), .A2(new_n459), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(G110), .B(G122), .Z(new_n505));
  NAND2_X1  g319(.A1(new_n261), .A2(new_n262), .ZN(new_n506));
  INV_X1    g320(.A(new_n210), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n418), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n463), .A3(G116), .ZN(new_n510));
  OAI211_X1 g324(.A(G113), .B(new_n510), .C1(new_n411), .C2(new_n509), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n415), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n248), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n505), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  INV_X1    g329(.A(new_n505), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n516), .C1(new_n263), .C2(new_n418), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(KEYINPUT6), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n192), .B(G125), .C1(new_n189), .C2(new_n193), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n519), .A2(KEYINPUT80), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(KEYINPUT80), .C1(G125), .C2(new_n237), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n244), .A2(G224), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT6), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n526), .B(new_n505), .C1(new_n508), .C2(new_n513), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n518), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n523), .B2(new_n524), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n520), .A2(new_n521), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n529), .A3(new_n522), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n248), .B2(new_n512), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n515), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n505), .B(KEYINPUT8), .Z(new_n538));
  NAND4_X1  g352(.A1(new_n230), .A2(new_n535), .A3(new_n415), .A4(new_n511), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(new_n517), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n528), .A2(new_n188), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G210), .B1(G237), .B2(G902), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT82), .Z(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n528), .A2(new_n188), .A3(new_n543), .A4(new_n541), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G214), .B1(G237), .B2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(KEYINPUT83), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n393), .A2(new_n504), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  NAND2_X1  g369(.A1(new_n438), .A2(new_n188), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n556), .A2(G472), .B1(new_n439), .B2(new_n438), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n496), .A2(KEYINPUT77), .A3(new_n497), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n557), .B(new_n279), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n503), .A2(new_n498), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(KEYINPUT92), .A3(new_n279), .A4(new_n557), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n565));
  INV_X1    g379(.A(new_n543), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n542), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n546), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n542), .B2(new_n566), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n548), .B(new_n392), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n379), .A2(new_n354), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT95), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n379), .A2(new_n573), .A3(new_n354), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n378), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT33), .B1(new_n378), .B2(KEYINPUT94), .ZN(new_n578));
  OAI211_X1 g392(.A(G478), .B(new_n188), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n350), .A2(new_n580), .A3(new_n352), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n570), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n562), .A2(new_n564), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT34), .B(G104), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G6));
  INV_X1    g399(.A(new_n385), .ZN(new_n586));
  INV_X1    g400(.A(new_n349), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n570), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n562), .A2(new_n564), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G107), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G9));
  NOR2_X1   g406(.A1(new_n489), .A2(KEYINPUT36), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n485), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n485), .A2(new_n594), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n597), .A2(new_n188), .A3(new_n462), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n496), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n393), .A2(new_n553), .A3(new_n557), .A4(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n601), .B(KEYINPUT37), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G110), .ZN(G12));
  AOI22_X1  g417(.A1(new_n441), .A2(new_n443), .B1(new_n458), .B2(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n274), .A2(new_n278), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n604), .A2(new_n605), .A3(new_n599), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n387), .B(KEYINPUT96), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(G900), .B2(new_n391), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n609), .B(KEYINPUT97), .Z(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n586), .A2(new_n587), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n548), .B1(new_n568), .B2(new_n569), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n606), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT99), .B(G128), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G30));
  XNOR2_X1  g433(.A(new_n547), .B(KEYINPUT100), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n610), .B(KEYINPUT39), .Z(new_n625));
  NAND2_X1  g439(.A1(new_n279), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT40), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n455), .A2(new_n425), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n450), .A2(new_n434), .A3(new_n426), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n444), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n350), .A2(new_n352), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(new_n548), .A3(new_n586), .A4(new_n636), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n624), .A2(new_n627), .A3(new_n600), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(new_n235), .ZN(G45));
  NAND4_X1  g453(.A1(new_n350), .A2(new_n580), .A3(new_n352), .A4(new_n611), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n606), .A2(new_n616), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G146), .ZN(G48));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n444), .A2(new_n459), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n260), .A2(new_n267), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n188), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(G469), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n278), .A3(new_n268), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n563), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n350), .A2(new_n352), .A3(new_n580), .ZN(new_n652));
  INV_X1    g466(.A(new_n569), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n546), .A3(new_n567), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n654), .A3(new_n548), .A4(new_n392), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n644), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n582), .A2(new_n504), .A3(KEYINPUT102), .A4(new_n650), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT41), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G113), .ZN(G15));
  NAND3_X1  g474(.A1(new_n589), .A2(new_n504), .A3(new_n650), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  NOR2_X1   g476(.A1(new_n615), .A2(new_n649), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n353), .A2(new_n385), .A3(new_n392), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n645), .A4(new_n600), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G119), .ZN(G21));
  NAND3_X1  g480(.A1(new_n586), .A2(new_n350), .A3(new_n352), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n570), .A2(new_n667), .ZN(new_n668));
  OR3_X1    g482(.A1(new_n496), .A2(KEYINPUT103), .A3(new_n497), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n428), .B(new_n437), .C1(new_n425), .C2(new_n453), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n556), .A2(G472), .B1(new_n439), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT103), .B1(new_n496), .B2(new_n497), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n668), .A2(new_n673), .A3(new_n650), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G122), .ZN(G24));
  NAND2_X1  g489(.A1(new_n641), .A2(KEYINPUT104), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n640), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n600), .A2(new_n671), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n663), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G125), .ZN(G27));
  INV_X1    g496(.A(new_n548), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n547), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n279), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n678), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n640), .A2(new_n677), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n504), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n685), .B1(new_n676), .B2(new_n678), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n669), .A2(new_n672), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n604), .A3(new_n690), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n222), .ZN(G33));
  NAND3_X1  g509(.A1(new_n614), .A2(new_n504), .A3(new_n686), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G134), .ZN(G36));
  AND2_X1   g511(.A1(new_n353), .A2(new_n580), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n699));
  OR3_X1    g513(.A1(new_n698), .A2(KEYINPUT106), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n557), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n699), .B1(new_n698), .B2(KEYINPUT106), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n600), .A4(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n684), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n256), .A2(new_n258), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n246), .B1(new_n709), .B2(new_n242), .ZN(new_n710));
  INV_X1    g524(.A(new_n269), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT45), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(G469), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n273), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n268), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n273), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n716), .A2(new_n722), .A3(new_n268), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n278), .A3(new_n625), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n705), .A2(new_n706), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n707), .A2(new_n708), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G137), .ZN(G39));
  NOR4_X1   g542(.A1(new_n563), .A2(new_n640), .A3(new_n683), .A4(new_n547), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n724), .B2(new_n278), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n724), .A2(new_n730), .A3(new_n278), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT47), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n733), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n604), .B(new_n729), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G140), .ZN(G42));
  OAI21_X1  g553(.A(new_n736), .B1(new_n735), .B2(new_n731), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n732), .A2(KEYINPUT47), .A3(new_n733), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n648), .A2(new_n268), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n740), .B(new_n741), .C1(new_n278), .C2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n700), .A2(new_n607), .A3(new_n702), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n673), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n684), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n548), .B1(new_n622), .B2(new_n623), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n744), .A2(new_n650), .A3(new_n673), .A4(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT50), .Z(new_n749));
  NAND2_X1  g563(.A1(new_n650), .A2(new_n684), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT117), .Z(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n635), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n563), .A3(new_n387), .A4(new_n753), .ZN(new_n754));
  OR3_X1    g568(.A1(new_n754), .A2(new_n636), .A3(new_n580), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n680), .A3(new_n744), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n746), .A2(new_n749), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n754), .A2(new_n581), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n386), .B(new_n761), .C1(new_n663), .C2(new_n745), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n760), .ZN(new_n764));
  INV_X1    g578(.A(new_n392), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n551), .B2(new_n552), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n636), .A2(new_n385), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n562), .A2(new_n564), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(new_n601), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n768), .B2(new_n601), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n562), .A2(new_n564), .A3(new_n766), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n554), .B1(new_n772), .B2(new_n581), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n599), .A2(new_n605), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n586), .A2(new_n349), .A3(new_n610), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n645), .A2(new_n775), .A3(new_n684), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n679), .A2(new_n680), .A3(new_n686), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n696), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n694), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n661), .A2(new_n674), .A3(new_n665), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n658), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT110), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n658), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n774), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n783), .A2(new_n786), .A3(new_n658), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n786), .B1(new_n783), .B2(new_n658), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(KEYINPUT113), .A3(new_n782), .A4(new_n774), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n606), .B(new_n616), .C1(new_n614), .C2(new_n641), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n279), .A2(new_n599), .A3(new_n611), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n615), .A2(new_n667), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n279), .A2(KEYINPUT114), .A3(new_n599), .A4(new_n611), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n635), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n681), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n795), .A2(new_n681), .A3(KEYINPUT52), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n790), .A2(new_n794), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n804), .A2(KEYINPUT115), .A3(new_n805), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n802), .A2(new_n811), .A3(new_n803), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n790), .A2(new_n794), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n808), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n784), .A2(new_n809), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n810), .A2(new_n816), .A3(new_n782), .A4(new_n812), .ZN(new_n817));
  INV_X1    g631(.A(new_n774), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(KEYINPUT54), .B(new_n819), .C1(new_n807), .C2(new_n809), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n815), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n808), .A2(new_n814), .A3(KEYINPUT116), .A4(KEYINPUT54), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n763), .A2(new_n764), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n692), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n752), .A2(new_n645), .A3(new_n825), .A4(new_n744), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT119), .Z(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT48), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n824), .A2(new_n828), .B1(G952), .B2(G953), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n692), .B1(KEYINPUT49), .B2(new_n742), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n548), .A3(new_n278), .A4(new_n698), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT109), .Z(new_n832));
  OR2_X1    g646(.A1(new_n742), .A2(KEYINPUT49), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n753), .A3(new_n624), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n834), .ZN(G75));
  NAND2_X1  g649(.A1(new_n518), .A2(new_n527), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n525), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT55), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n819), .B1(new_n807), .B2(new_n809), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n188), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(G210), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n244), .A2(G952), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n842), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n840), .B2(new_n544), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(G51));
  NAND2_X1  g661(.A1(new_n273), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n807), .A2(new_n809), .ZN(new_n850));
  INV_X1    g664(.A(new_n819), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n848), .B1(new_n852), .B2(new_n820), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n273), .A2(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n646), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n839), .A2(new_n188), .A3(new_n715), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n844), .B1(new_n855), .B2(new_n856), .ZN(G54));
  NAND3_X1  g671(.A1(new_n840), .A2(KEYINPUT58), .A3(G475), .ZN(new_n858));
  INV_X1    g672(.A(new_n344), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n858), .A2(KEYINPUT120), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n844), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n858), .B2(new_n859), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT120), .B1(new_n858), .B2(new_n859), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(G60));
  OR2_X1    g678(.A1(new_n577), .A2(new_n578), .ZN(new_n865));
  NAND2_X1  g679(.A1(G478), .A2(G902), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT59), .Z(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n865), .B(new_n868), .C1(new_n852), .C2(new_n820), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n869), .A2(new_n861), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n822), .B2(new_n823), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n870), .B(KEYINPUT121), .C1(new_n865), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n821), .B1(new_n839), .B2(new_n849), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n808), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n823), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n865), .B1(new_n876), .B2(new_n868), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n869), .A2(new_n861), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n879), .ZN(G63));
  NAND2_X1  g694(.A1(new_n850), .A2(new_n851), .ZN(new_n881));
  NAND2_X1  g695(.A1(G217), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT60), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n490), .A2(new_n491), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n844), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n881), .A2(new_n597), .A3(new_n884), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n839), .A2(new_n883), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(KEYINPUT122), .A3(new_n597), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT122), .B1(new_n891), .B2(new_n597), .ZN(new_n899));
  INV_X1    g713(.A(new_n597), .ZN(new_n900));
  NOR4_X1   g714(.A1(new_n839), .A2(new_n889), .A3(new_n900), .A4(new_n883), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n894), .A3(new_n895), .A4(new_n887), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n898), .A2(new_n903), .ZN(G66));
  AOI21_X1  g718(.A(new_n244), .B1(new_n389), .B2(G224), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n793), .A2(new_n774), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n907), .B2(new_n244), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n836), .B1(G898), .B2(new_n244), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(G69));
  AOI21_X1  g724(.A(new_n244), .B1(G227), .B2(G900), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n403), .A2(new_n409), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n328), .A2(new_n330), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT124), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n912), .B(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n244), .A2(G900), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n725), .A2(new_n645), .A3(new_n825), .A4(new_n799), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n795), .A2(new_n681), .ZN(new_n918));
  INV_X1    g732(.A(new_n696), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n694), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n738), .A2(new_n727), .A3(new_n917), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n921), .B2(new_n244), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n924), .B(new_n916), .C1(new_n921), .C2(new_n244), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n915), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n911), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n638), .A2(new_n918), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n581), .B1(new_n636), .B2(new_n385), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n504), .A2(new_n931), .A3(new_n686), .A4(new_n625), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n738), .A2(new_n930), .A3(new_n727), .A4(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(new_n244), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(new_n915), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n926), .B(new_n935), .C1(new_n927), .C2(new_n911), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G72));
  NAND2_X1  g753(.A1(G472), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT63), .Z(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n921), .B2(new_n907), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n844), .B1(new_n942), .B2(new_n456), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n933), .B2(new_n907), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n425), .A3(new_n455), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n628), .A2(new_n941), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n808), .A2(new_n457), .A3(new_n814), .A4(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G57));
endmodule


