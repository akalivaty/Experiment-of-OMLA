//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G134gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n204), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g017(.A(G148gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(G141gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT70), .B(G141gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n214), .B1(new_n223), .B2(new_n215), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n218), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n212), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G225gat), .A2(G233gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n212), .A2(new_n225), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OR3_X1    g033(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n235));
  OAI211_X1 g034(.A(KEYINPUT72), .B(new_n232), .C1(new_n212), .C2(new_n225), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n212), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n240), .A2(new_n227), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n237), .A2(KEYINPUT73), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT73), .B1(new_n237), .B2(new_n241), .ZN(new_n243));
  OAI211_X1 g042(.A(KEYINPUT5), .B(new_n229), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n231), .A2(new_n232), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(new_n240), .C1(KEYINPUT4), .C2(new_n231), .ZN(new_n246));
  OR3_X1    g045(.A1(new_n246), .A2(KEYINPUT5), .A3(new_n228), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G1gat), .B(G29gat), .Z(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G57gat), .B(G85gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n255));
  INV_X1    g054(.A(new_n253), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n244), .A2(new_n256), .A3(new_n247), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n253), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G8gat), .ZN(new_n263));
  INV_X1    g062(.A(G36gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(KEYINPUT64), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(KEYINPUT27), .B2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(new_n267), .C1(new_n266), .C2(KEYINPUT64), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT27), .B(G183gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT28), .A3(new_n267), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT26), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n276), .B(new_n282), .C1(new_n280), .C2(new_n279), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n267), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT23), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n281), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  OR2_X1    g088(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n290), .A2(G190gat), .A3(new_n291), .ZN(new_n292));
  OR3_X1    g091(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n288), .B2(new_n292), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n283), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT68), .B(KEYINPUT29), .Z(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n309), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n308), .B(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n297), .B1(new_n296), .B2(KEYINPUT29), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n265), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n317), .B2(new_n316), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n311), .A2(KEYINPUT30), .A3(new_n315), .A4(new_n265), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n260), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT34), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n283), .A2(new_n295), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n212), .ZN(new_n325));
  INV_X1    g124(.A(G227gat), .ZN(new_n326));
  INV_X1    g125(.A(G233gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n212), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n283), .A2(new_n295), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n323), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  INV_X1    g137(.A(new_n331), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n330), .B1(new_n283), .B2(new_n295), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n328), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT66), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n331), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT66), .B1(new_n344), .B2(new_n328), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n338), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G15gat), .B(G43gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND3_X1  g148(.A1(new_n337), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n341), .A2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(KEYINPUT66), .A3(new_n328), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT33), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n349), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n335), .B(new_n336), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT32), .B1(new_n343), .B2(new_n345), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n350), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n350), .B2(new_n355), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT82), .B(G22gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n310), .A2(new_n300), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n225), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n300), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n238), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n310), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n372), .B(KEYINPUT78), .Z(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n313), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n364), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n225), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n372), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n370), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n376), .A2(new_n377), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n364), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n372), .B1(new_n388), .B2(new_n225), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT81), .B1(new_n389), .B2(new_n370), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n361), .B(new_n374), .C1(new_n385), .C2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT76), .B(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT75), .B(KEYINPUT31), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G22gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n373), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n367), .B2(new_n370), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n389), .A2(KEYINPUT81), .A3(new_n370), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n391), .B(new_n396), .C1(new_n397), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n396), .B(KEYINPUT77), .Z(new_n405));
  OAI21_X1  g204(.A(new_n374), .B1(new_n385), .B2(new_n390), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n360), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n391), .ZN(new_n408));
  OAI22_X1  g207(.A1(new_n358), .A2(new_n359), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT35), .B1(new_n322), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n350), .A2(new_n355), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n356), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n350), .A2(new_n355), .A3(new_n357), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n402), .B(new_n360), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n403), .B1(new_n417), .B2(new_n405), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n260), .A3(new_n418), .A4(new_n321), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT87), .B1(new_n419), .B2(KEYINPUT35), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n260), .A2(new_n321), .ZN(new_n421));
  INV_X1    g220(.A(new_n409), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT35), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(KEYINPUT88), .A3(KEYINPUT35), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n412), .A2(new_n420), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n319), .A2(new_n320), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT40), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n248), .B2(new_n253), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n246), .A2(new_n228), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n432), .A2(KEYINPUT39), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n432), .B(KEYINPUT39), .C1(new_n228), .C2(new_n226), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n433), .A2(new_n434), .A3(new_n256), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n436), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n428), .A2(new_n431), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n316), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n441), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n315), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n316), .A2(KEYINPUT37), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT38), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n302), .A2(new_n313), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n299), .A2(new_n310), .A3(new_n314), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT84), .A4(KEYINPUT37), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n451), .A2(new_n265), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT38), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(KEYINPUT37), .A3(new_n450), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n445), .A2(new_n452), .A3(new_n453), .A4(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n448), .A2(new_n259), .A3(new_n457), .A4(new_n258), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n265), .B1(new_n316), .B2(new_n453), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n418), .B(new_n439), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n418), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n322), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n416), .B(KEYINPUT36), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n427), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(G15gat), .A2(G22gat), .ZN(new_n466));
  INV_X1    g265(.A(G1gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(G15gat), .A2(G22gat), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(KEYINPUT16), .ZN(new_n470));
  AND2_X1   g269(.A1(G15gat), .A2(G22gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(G15gat), .A2(G22gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G8gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n466), .A2(new_n468), .B1(KEYINPUT16), .B2(new_n467), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n471), .A2(new_n472), .A3(G1gat), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT91), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT92), .B(G8gat), .Z(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT93), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n474), .B2(KEYINPUT91), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT93), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n481), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n476), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G71gat), .A2(G78gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT96), .ZN(new_n493));
  INV_X1    g292(.A(G64gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G57gat), .ZN(new_n495));
  INV_X1    g294(.A(G57gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G64gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n490), .A2(new_n500), .A3(new_n491), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n493), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n490), .B(new_n503), .C1(new_n504), .C2(new_n491), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT21), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G183gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n266), .A3(new_n507), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n514));
  INV_X1    g313(.A(G231gat), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n327), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n511), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT97), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(new_n327), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n512), .ZN(new_n520));
  XNOR2_X1  g319(.A(G127gat), .B(G155gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n305), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n516), .B2(new_n520), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n506), .A2(KEYINPUT21), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n527), .B(new_n528), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n520), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n533), .B2(new_n524), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n264), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT89), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT15), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT15), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  INV_X1    g348(.A(G43gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(G50gat), .ZN(new_n551));
  INV_X1    g350(.A(G50gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G43gat), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT90), .B(new_n549), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n540), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n548), .A2(new_n554), .A3(new_n555), .A4(new_n542), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n546), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n563), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n577), .A2(new_n572), .A3(new_n566), .A4(new_n570), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n566), .A2(new_n570), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT99), .A3(new_n572), .A4(new_n577), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(KEYINPUT100), .A3(new_n573), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n576), .A2(new_n580), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n561), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT98), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n586), .A2(new_n557), .B1(KEYINPUT41), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n589), .A2(KEYINPUT41), .ZN(new_n595));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n591), .A2(new_n592), .ZN(new_n599));
  OR3_X1    g398(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n594), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n535), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n465), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT10), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n584), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n574), .A2(KEYINPUT101), .A3(new_n578), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n571), .A2(new_n608), .A3(new_n573), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n506), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n584), .B2(new_n506), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT102), .B(KEYINPUT10), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n606), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT105), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n580), .A2(new_n582), .ZN(new_n619));
  INV_X1    g418(.A(new_n506), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n571), .A2(KEYINPUT100), .A3(new_n573), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT100), .B1(new_n571), .B2(new_n573), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n612), .B1(new_n624), .B2(new_n610), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n618), .B(new_n615), .C1(new_n625), .C2(new_n606), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n611), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n616), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n278), .ZN(new_n631));
  INV_X1    g430(.A(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT104), .Z(new_n634));
  NOR2_X1   g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n625), .A2(KEYINPUT103), .A3(new_n606), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n611), .A2(new_n613), .ZN(new_n638));
  INV_X1    g437(.A(new_n606), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n615), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n628), .A2(new_n616), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n561), .A2(new_n489), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n487), .B1(new_n486), .B2(new_n481), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n480), .B1(new_n469), .B2(new_n473), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n466), .A2(new_n468), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT91), .B1(new_n651), .B2(new_n470), .ZN(new_n652));
  NOR4_X1   g451(.A1(new_n650), .A2(new_n652), .A3(KEYINPUT93), .A4(new_n482), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n475), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n557), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(new_n648), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(KEYINPUT18), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT95), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT11), .B(G169gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G197gat), .ZN(new_n663));
  XOR2_X1   g462(.A(G113gat), .B(G141gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n648), .B(KEYINPUT13), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n655), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n654), .A2(new_n557), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n647), .A2(new_n655), .A3(KEYINPUT18), .A4(new_n648), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n660), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n673), .A3(new_n674), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n661), .A3(new_n667), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n646), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n604), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n260), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n258), .A2(KEYINPUT106), .A3(new_n259), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g489(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n691));
  OR2_X1    g490(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n683), .A2(new_n428), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n683), .ZN(new_n696));
  OAI21_X1  g495(.A(G8gat), .B1(new_n696), .B2(new_n321), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(G1325gat));
  AOI21_X1  g498(.A(G15gat), .B1(new_n683), .B2(new_n416), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT36), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n416), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G15gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT107), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n700), .B1(new_n683), .B2(new_n704), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n683), .A2(new_n461), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NAND2_X1  g507(.A1(new_n465), .A2(new_n602), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n531), .A2(new_n534), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n682), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n537), .A3(new_n688), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n602), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n427), .B2(new_n464), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT44), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n715), .A2(new_n681), .A3(new_n535), .A4(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n687), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n720), .ZN(G1328gat));
  AND3_X1   g520(.A1(new_n711), .A2(new_n264), .A3(new_n428), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n719), .B2(new_n321), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n724), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(G1329gat));
  OAI21_X1  g527(.A(G43gat), .B1(new_n719), .B2(new_n463), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n550), .A3(new_n416), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  OAI21_X1  g533(.A(G50gat), .B1(new_n719), .B2(new_n418), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n711), .A2(new_n552), .A3(new_n461), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n735), .B(new_n738), .C1(new_n736), .C2(KEYINPUT48), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1331gat));
  NOR2_X1   g542(.A1(new_n645), .A2(new_n679), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n465), .A2(new_n603), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n687), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n496), .ZN(G1332gat));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n321), .ZN(new_n748));
  NOR2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  AND2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n748), .B2(new_n749), .ZN(G1333gat));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  INV_X1    g552(.A(G71gat), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n745), .A2(new_n754), .A3(new_n463), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(new_n416), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n416), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n754), .B1(new_n745), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n756), .A2(new_n757), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n757), .B1(new_n756), .B2(new_n763), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n753), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n766), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(KEYINPUT50), .A3(new_n764), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1334gat));
  NOR2_X1   g569(.A1(new_n745), .A2(new_n418), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(G78gat), .Z(G1335gat));
  AOI21_X1  g571(.A(new_n710), .B1(new_n709), .B2(new_n714), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(new_n718), .A3(new_n744), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n774), .A2(new_n567), .A3(new_n687), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n465), .A2(new_n680), .A3(new_n535), .A4(new_n602), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n717), .A2(KEYINPUT51), .A3(new_n680), .A4(new_n535), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AOI211_X1 g580(.A(new_n710), .B(new_n716), .C1(new_n427), .C2(new_n464), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n680), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n781), .A2(new_n688), .A3(new_n646), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n775), .B1(new_n567), .B2(new_n784), .ZN(G1336gat));
  NAND3_X1  g584(.A1(new_n778), .A2(KEYINPUT113), .A3(new_n780), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n321), .A2(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n776), .A2(new_n788), .A3(new_n777), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n786), .A2(new_n646), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n428), .A3(new_n718), .A4(new_n744), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n781), .A2(new_n646), .A3(new_n783), .A4(new_n787), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  OAI21_X1  g596(.A(G92gat), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n535), .B1(new_n717), .B2(KEYINPUT44), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n714), .B(new_n716), .C1(new_n427), .C2(new_n464), .ZN(new_n800));
  INV_X1    g599(.A(new_n744), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT114), .B1(new_n802), .B2(new_n428), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n795), .B(new_n796), .C1(new_n798), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n794), .A2(new_n804), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n774), .B2(new_n463), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n758), .A2(G99gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n781), .A2(new_n646), .A3(new_n783), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n808), .A3(KEYINPUT115), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  OAI21_X1  g612(.A(G106gat), .B1(new_n774), .B2(new_n418), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n418), .A2(G106gat), .A3(new_n645), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n781), .A2(new_n783), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n786), .A2(new_n789), .A3(new_n816), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n815), .ZN(G1339gat));
  NAND2_X1  g620(.A1(new_n614), .A2(new_n616), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n642), .B1(new_n627), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n644), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n825), .A3(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n823), .A2(new_n825), .A3(new_n831), .A4(KEYINPUT55), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n828), .A2(new_n830), .A3(new_n679), .A4(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n671), .A2(new_n672), .A3(new_n670), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n648), .B1(new_n647), .B2(new_n655), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n665), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n675), .A2(new_n666), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n836), .B(new_n837), .C1(new_n635), .C2(new_n644), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n602), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n828), .A2(new_n830), .A3(new_n832), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n602), .A2(new_n836), .A3(new_n837), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n535), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n710), .A2(new_n680), .A3(new_n645), .A4(new_n716), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n685), .A2(new_n686), .A3(new_n321), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n409), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n679), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n646), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n848), .A2(new_n535), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(new_n208), .ZN(G1342gat));
  NOR2_X1   g654(.A1(new_n848), .A2(new_n716), .ZN(new_n856));
  INV_X1    g655(.A(G134gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n859), .B(new_n860), .C1(new_n857), .C2(new_n856), .ZN(G1343gat));
  AOI21_X1  g660(.A(new_n418), .B1(new_n843), .B2(new_n844), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n702), .A2(new_n846), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G141gat), .A3(new_n680), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT57), .B(new_n418), .C1(new_n843), .C2(new_n844), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n869), .A2(new_n680), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n866), .B1(new_n221), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n463), .A2(new_n688), .A3(new_n321), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n845), .A2(new_n461), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n867), .ZN(new_n876));
  INV_X1    g675(.A(new_n870), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n870), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n679), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n221), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n865), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n872), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT119), .B(new_n872), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1344gat));
  INV_X1    g687(.A(new_n864), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n219), .A3(new_n646), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n867), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(KEYINPUT57), .B2(new_n875), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n646), .A3(new_n863), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n219), .B1(new_n894), .B2(KEYINPUT120), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n878), .A2(new_n879), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n891), .B1(new_n898), .B2(new_n645), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n219), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n890), .B1(new_n897), .B2(new_n900), .ZN(G1345gat));
  AOI21_X1  g700(.A(G155gat), .B1(new_n889), .B2(new_n710), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n898), .A2(new_n535), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g703(.A(G162gat), .B1(new_n889), .B2(new_n602), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n898), .A2(new_n716), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(G162gat), .ZN(G1347gat));
  NAND2_X1  g706(.A1(new_n845), .A2(new_n687), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n845), .A2(new_n910), .A3(new_n687), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n409), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n428), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n277), .A3(new_n679), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n759), .A2(new_n418), .A3(new_n761), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n845), .A2(new_n916), .A3(new_n687), .A4(new_n428), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n680), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(G1348gat));
  NOR3_X1   g718(.A1(new_n917), .A2(new_n278), .A3(new_n645), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n914), .A2(new_n646), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n278), .ZN(G1349gat));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n710), .A3(new_n274), .ZN(new_n923));
  OAI21_X1  g722(.A(G183gat), .B1(new_n917), .B2(new_n535), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(G190gat), .C1(new_n917), .C2(new_n716), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n917), .A2(new_n716), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G190gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n934), .B2(KEYINPUT61), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT123), .B(new_n927), .C1(new_n933), .C2(G190gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n931), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n716), .A2(G190gat), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT122), .B1(new_n913), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n912), .A2(new_n941), .A3(new_n428), .A4(new_n938), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT125), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n940), .A2(new_n942), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n935), .A2(new_n936), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n945), .B(new_n946), .C1(new_n947), .C2(new_n931), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(new_n948), .ZN(G1351gat));
  NAND3_X1  g748(.A1(new_n463), .A2(new_n687), .A3(new_n428), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n893), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(new_n680), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(G197gat), .A3(new_n955), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n321), .B(new_n702), .C1(new_n909), .C2(new_n911), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n461), .ZN(new_n958));
  OR3_X1    g757(.A1(new_n958), .A2(G197gat), .A3(new_n680), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n956), .A2(new_n959), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n646), .A2(new_n632), .ZN(new_n961));
  OR3_X1    g760(.A1(new_n958), .A2(KEYINPUT62), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n958), .B2(new_n961), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n951), .A2(new_n893), .A3(new_n646), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n962), .B(new_n963), .C1(new_n632), .C2(new_n964), .ZN(G1353gat));
  NAND4_X1  g764(.A1(new_n957), .A2(new_n305), .A3(new_n710), .A4(new_n461), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n893), .A2(new_n710), .A3(new_n951), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  OAI21_X1  g769(.A(G218gat), .B1(new_n952), .B2(new_n716), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n602), .A2(new_n306), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n958), .B2(new_n972), .ZN(G1355gat));
endmodule


