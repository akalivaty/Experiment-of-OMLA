//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n191), .A2(G146), .A3(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT67), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n200), .A3(G128), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n201), .A2(KEYINPUT73), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n201), .B(KEYINPUT73), .C1(new_n197), .C2(G128), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT24), .B(G110), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(G119), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(KEYINPUT23), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n198), .A2(new_n200), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(KEYINPUT74), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G110), .ZN(new_n216));
  OAI221_X1 g030(.A(new_n196), .B1(new_n204), .B2(new_n205), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n216), .A3(new_n214), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n191), .A2(G146), .A3(new_n192), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT75), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  AOI211_X1 g042(.A(new_n228), .B(new_n225), .C1(new_n218), .C2(new_n219), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n217), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT77), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G137), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT76), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT76), .B(new_n217), .C1(new_n227), .C2(new_n229), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n235), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G234), .ZN(new_n243));
  OAI21_X1  g057(.A(G217), .B1(new_n243), .B2(G902), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT78), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n248));
  INV_X1    g062(.A(new_n246), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n248), .B(new_n249), .C1(new_n250), .C2(new_n236), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(new_n245), .C1(new_n250), .C2(new_n236), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n244), .B(KEYINPUT72), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n245), .B1(new_n250), .B2(new_n236), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(KEYINPUT25), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n264));
  OAI211_X1 g078(.A(G134), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n262), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n265), .A2(new_n266), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(new_n264), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n273), .B2(new_n262), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT80), .ZN(new_n276));
  INV_X1    g090(.A(G104), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT3), .B1(new_n277), .B2(G107), .ZN(new_n278));
  AOI21_X1  g092(.A(G101), .B1(new_n277), .B2(G107), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n280));
  INV_X1    g094(.A(G107), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G104), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G101), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(G107), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(G104), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n276), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n223), .A2(G143), .ZN(new_n289));
  INV_X1    g103(.A(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G146), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(KEYINPUT1), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(G128), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n289), .B(new_n291), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(new_n286), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G101), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT80), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n294), .A2(new_n298), .A3(new_n295), .A4(new_n299), .ZN(new_n302));
  AOI221_X4 g116(.A(new_n260), .B1(new_n271), .B2(new_n275), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n275), .A2(new_n271), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT12), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT0), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n211), .A3(KEYINPUT64), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(KEYINPUT0), .B2(G128), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n292), .A2(new_n308), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G143), .B(G146), .ZN(new_n314));
  INV_X1    g128(.A(new_n308), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT65), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n310), .A2(new_n312), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(KEYINPUT65), .A3(new_n292), .A4(new_n308), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n278), .A2(new_n282), .A3(new_n285), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G101), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT4), .A3(new_n299), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n324), .A3(G101), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n294), .A2(new_n295), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT80), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT80), .B1(new_n298), .B2(new_n299), .ZN(new_n329));
  OAI211_X1 g143(.A(KEYINPUT10), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n305), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT10), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n302), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n326), .A2(new_n330), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n231), .A2(G227), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n259), .B1(new_n307), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n304), .A2(new_n305), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n260), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n304), .A2(KEYINPUT12), .A3(new_n305), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n334), .A2(new_n338), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT81), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n323), .A2(new_n325), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n347), .A2(new_n320), .B1(new_n332), .B2(new_n302), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n331), .B1(new_n348), .B2(new_n330), .ZN(new_n349));
  INV_X1    g163(.A(new_n334), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n337), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n340), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n245), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n245), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n334), .B1(new_n303), .B2(new_n306), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n337), .B(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n330), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n305), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n356), .A2(new_n357), .B1(new_n359), .B2(new_n345), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n355), .B1(new_n360), .B2(G469), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT9), .B(G234), .ZN(new_n363));
  OAI21_X1  g177(.A(G221), .B1(new_n363), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(KEYINPUT20), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(KEYINPUT20), .ZN(new_n367));
  NOR2_X1   g181(.A1(G237), .A2(G953), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G143), .A3(G214), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(G143), .B1(new_n368), .B2(G214), .ZN(new_n371));
  OAI21_X1  g185(.A(G131), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT17), .ZN(new_n373));
  INV_X1    g187(.A(G237), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n231), .A3(G214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n290), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n266), .A3(new_n369), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n266), .B1(new_n376), .B2(new_n369), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n379), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT89), .B1(new_n379), .B2(KEYINPUT17), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n195), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n277), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT18), .B(G131), .C1(new_n370), .C2(new_n371), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n188), .A2(new_n190), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n224), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n376), .A2(new_n369), .A3(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n385), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n382), .A2(new_n384), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT19), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT19), .B1(new_n188), .B2(new_n190), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n223), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT19), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n222), .A2(KEYINPUT19), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT87), .A3(new_n223), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n193), .B1(new_n372), .B2(new_n377), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n391), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n384), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n396), .A2(new_n397), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n402), .B2(new_n223), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n392), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT88), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n393), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(G475), .A2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n366), .B(new_n367), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n382), .A2(new_n384), .A3(new_n392), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n407), .A3(new_n392), .ZN(new_n419));
  INV_X1    g233(.A(new_n384), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n406), .A2(new_n407), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(new_n365), .A3(KEYINPUT20), .A4(new_n415), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n384), .B1(new_n382), .B2(new_n392), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n245), .B1(new_n393), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G475), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n417), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT93), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT14), .B1(new_n433), .B2(G116), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G116), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G122), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(G116), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n438), .B2(KEYINPUT14), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n281), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n438), .A2(new_n441), .A3(new_n281), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n290), .A2(G128), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n211), .A2(G143), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n267), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n267), .B1(new_n446), .B2(new_n447), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT92), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n438), .A2(new_n441), .A3(new_n281), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n281), .B1(new_n438), .B2(new_n441), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT13), .B1(new_n290), .B2(G128), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n290), .A2(G128), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n290), .A2(KEYINPUT13), .A3(G128), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n267), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n446), .A2(new_n447), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G134), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n453), .B1(new_n464), .B2(new_n448), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n442), .B1(new_n436), .B2(new_n439), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n465), .B(new_n466), .C1(new_n281), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n452), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G217), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n363), .A2(new_n470), .A3(G953), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n452), .A2(new_n462), .A3(new_n468), .A4(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n432), .B1(new_n475), .B2(new_n245), .ZN(new_n476));
  AOI211_X1 g290(.A(KEYINPUT93), .B(G902), .C1(new_n473), .C2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n431), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n465), .B1(new_n281), .B2(new_n467), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n461), .B1(new_n479), .B2(KEYINPUT92), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n471), .B1(new_n480), .B2(new_n468), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n468), .A2(new_n452), .A3(new_n462), .A4(new_n471), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n245), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n431), .B1(new_n483), .B2(KEYINPUT93), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n231), .A2(G952), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(G234), .B2(G237), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT21), .B(G898), .Z(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT94), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n245), .B(new_n231), .C1(G234), .C2(G237), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT95), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n478), .A2(new_n485), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n362), .A2(new_n364), .A3(new_n429), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G214), .B1(G237), .B2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n198), .A2(new_n200), .A3(G116), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n437), .A2(G119), .ZN(new_n498));
  INV_X1    g312(.A(G113), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT2), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT2), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G113), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT68), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n497), .A2(new_n503), .A3(new_n506), .A4(new_n498), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT82), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(KEYINPUT5), .A3(new_n498), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT82), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT5), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n207), .A2(new_n511), .A3(new_n512), .A4(G116), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n509), .A2(new_n510), .A3(G113), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n328), .A2(new_n329), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n497), .A2(new_n498), .ZN(new_n517));
  INV_X1    g331(.A(new_n503), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n505), .A2(new_n507), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n323), .A2(new_n325), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n515), .A2(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G110), .B(G122), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT83), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n347), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT83), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n508), .B(new_n514), .C1(new_n329), .C2(new_n328), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n522), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n522), .B1(new_n527), .B2(new_n529), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n521), .A2(new_n533), .A3(new_n523), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n317), .A2(new_n319), .A3(G125), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n296), .A2(new_n189), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n231), .A2(G224), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n535), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n538), .B2(KEYINPUT86), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n540), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n538), .B(new_n539), .C1(KEYINPUT86), .C2(new_n545), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n524), .B2(new_n530), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n522), .B(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n508), .A2(new_n514), .B1(new_n299), .B2(new_n298), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n529), .B1(new_n553), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n544), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n544), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n496), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n495), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n271), .A2(new_n275), .B1(new_n317), .B2(new_n319), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n269), .A2(new_n268), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G131), .ZN(new_n566));
  AND4_X1   g380(.A1(new_n271), .A2(new_n295), .A3(new_n294), .A4(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n564), .A2(new_n567), .A3(KEYINPUT30), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n305), .A2(new_n320), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n327), .A2(new_n271), .A3(new_n566), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n526), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n368), .A2(G210), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n519), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n570), .A2(new_n519), .A3(new_n571), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT30), .B1(new_n564), .B2(new_n567), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n570), .A2(new_n569), .A3(new_n571), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n586), .B2(new_n526), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT31), .A3(new_n578), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT28), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n526), .B1(new_n564), .B2(new_n567), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(new_n579), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n564), .A2(new_n567), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT28), .B1(new_n592), .B2(new_n519), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT70), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n519), .B1(new_n570), .B2(new_n571), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT28), .B1(new_n583), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT70), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n578), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n582), .A2(new_n588), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(G472), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT32), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n582), .A2(new_n588), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n579), .A2(new_n589), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n597), .B1(new_n596), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n591), .A2(KEYINPUT70), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT32), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n602), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT29), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n519), .B1(new_n584), .B2(new_n585), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n600), .B1(new_n615), .B2(new_n583), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n614), .B(new_n616), .C1(new_n599), .C2(new_n600), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT71), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n590), .B2(new_n579), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n595), .A2(KEYINPUT71), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT28), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n621), .A2(KEYINPUT29), .A3(new_n578), .A4(new_n606), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(new_n245), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n258), .A2(new_n563), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n562), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n559), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n542), .B(new_n536), .C1(new_n531), .C2(new_n534), .ZN(new_n631));
  INV_X1    g445(.A(new_n549), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n531), .A2(new_n557), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n245), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n630), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n544), .A2(new_n558), .A3(new_n559), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(KEYINPUT96), .A3(new_n496), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n430), .A2(G902), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(KEYINPUT97), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(KEYINPUT97), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n642), .B(new_n643), .C1(new_n473), .C2(new_n474), .ZN(new_n644));
  AND4_X1   g458(.A1(KEYINPUT97), .A2(new_n473), .A3(new_n641), .A4(new_n474), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n483), .A2(new_n430), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n428), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n639), .A2(new_n493), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n601), .B2(G902), .ZN(new_n651));
  INV_X1    g465(.A(new_n364), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n354), .B2(new_n361), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n610), .A2(new_n602), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n258), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  AOI21_X1  g473(.A(KEYINPUT98), .B1(new_n417), .B2(new_n424), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n478), .A2(new_n485), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n417), .A2(new_n424), .A3(KEYINPUT98), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n661), .A2(new_n427), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n639), .A2(new_n665), .A3(new_n493), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n656), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n281), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  NAND2_X1  g484(.A1(new_n651), .A2(new_n654), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n256), .A2(KEYINPUT25), .ZN(new_n673));
  INV_X1    g487(.A(new_n255), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n254), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT100), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n240), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n249), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n563), .A2(new_n672), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  AOI22_X1  g497(.A1(new_n604), .A2(new_n612), .B1(new_n623), .B2(G472), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n257), .A2(new_n254), .B1(new_n249), .B2(new_n678), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n491), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n487), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n664), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n686), .A2(new_n639), .A3(new_n653), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XNOR2_X1  g508(.A(new_n637), .B(KEYINPUT101), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n690), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n653), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT40), .Z(new_n701));
  NOR2_X1   g515(.A1(new_n619), .A2(new_n620), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n580), .B1(new_n702), .B2(new_n578), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n245), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n613), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n496), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n428), .A2(new_n662), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n707), .A2(new_n708), .A3(new_n680), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n698), .A2(new_n701), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n428), .A2(new_n648), .A3(new_n690), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n686), .A2(new_n639), .A3(new_n653), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  NAND2_X1  g530(.A1(new_n258), .A2(new_n625), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n352), .A2(new_n245), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n354), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(KEYINPUT103), .A3(G469), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT104), .B1(new_n723), .B2(new_n364), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n725), .B(new_n652), .C1(new_n721), .C2(new_n722), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n717), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n650), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  AND2_X1   g545(.A1(new_n247), .A2(new_n251), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n675), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n684), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n354), .A2(new_n720), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n353), .B1(new_n352), .B2(new_n245), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n722), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n364), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n725), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n652), .B1(new_n721), .B2(new_n722), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n734), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(new_n666), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT105), .B(G116), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G18));
  INV_X1    g560(.A(new_n493), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n428), .A2(new_n662), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n686), .A2(new_n639), .A3(new_n748), .A4(new_n741), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  AOI21_X1  g564(.A(new_n709), .B1(new_n629), .B2(new_n638), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n493), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n724), .A2(new_n726), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT107), .B1(new_n732), .B2(new_n675), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n258), .A2(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT31), .B1(new_n587), .B2(new_n578), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n615), .A2(new_n581), .A3(new_n600), .A4(new_n583), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n578), .B1(new_n621), .B2(new_n606), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n602), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(G902), .B1(new_n605), .B2(new_n609), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT106), .B(G472), .Z(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n752), .A2(new_n753), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  AOI21_X1  g583(.A(new_n766), .B1(new_n675), .B2(new_n679), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n639), .A2(new_n714), .A3(new_n770), .A4(new_n741), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G125), .ZN(G27));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n613), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n604), .A2(KEYINPUT108), .A3(new_n612), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n624), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n653), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n635), .A2(new_n496), .A3(new_n636), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n713), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n732), .A2(KEYINPUT107), .A3(new_n675), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n776), .B(new_n780), .C1(new_n754), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n777), .A2(new_n778), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n258), .A2(new_n625), .A3(new_n783), .A4(new_n714), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n779), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NAND4_X1  g601(.A1(new_n258), .A2(new_n692), .A3(new_n625), .A4(new_n783), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT109), .B(G134), .Z(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G36));
  AOI21_X1  g604(.A(new_n428), .B1(new_n647), .B2(new_n646), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT43), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n792), .A2(new_n671), .A3(new_n680), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n778), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(KEYINPUT112), .A3(KEYINPUT44), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n360), .A2(KEYINPUT45), .ZN(new_n804));
  OAI21_X1  g618(.A(G469), .B1(new_n360), .B2(KEYINPUT45), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n353), .B2(new_n245), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT46), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n807), .A2(KEYINPUT110), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT110), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n354), .A3(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n811), .A2(KEYINPUT111), .B1(new_n808), .B2(new_n807), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n809), .A2(new_n813), .A3(new_n354), .A4(new_n810), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n652), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n802), .A2(new_n699), .A3(new_n803), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  NOR4_X1   g631(.A1(new_n258), .A2(new_n625), .A3(new_n713), .A4(new_n778), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n815), .A2(KEYINPUT47), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n815), .A2(KEYINPUT47), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  NAND2_X1  g636(.A1(new_n741), .A2(new_n797), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n823), .A2(new_n706), .A3(new_n733), .A4(new_n689), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n429), .A3(new_n647), .A4(new_n646), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n680), .A2(new_n767), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n792), .A2(new_n487), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(new_n823), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n697), .A2(new_n708), .A3(new_n741), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n767), .B1(new_n781), .B2(new_n754), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n827), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(KEYINPUT50), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n830), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n830), .B2(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n829), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n723), .A2(new_n652), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n819), .A2(new_n820), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n797), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT51), .B(new_n838), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT96), .B1(new_n637), .B2(new_n496), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n628), .B(new_n708), .C1(new_n635), .C2(new_n636), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n741), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n833), .A2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n486), .B(new_n850), .C1(new_n649), .C2(new_n824), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n757), .A2(new_n776), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n827), .A2(new_n823), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT48), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT121), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n855), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n845), .B(new_n846), .C1(new_n856), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n483), .A2(KEYINPUT93), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n475), .A2(new_n432), .A3(new_n245), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n484), .B1(new_n864), .B2(new_n431), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n428), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n649), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n496), .B(new_n493), .C1(new_n560), .C2(new_n561), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n258), .A3(new_n655), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n626), .A3(new_n681), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n782), .B2(new_n785), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n625), .A2(new_n680), .A3(new_n748), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n849), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n727), .B2(new_n728), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n875), .A3(new_n744), .A4(new_n768), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n690), .A2(KEYINPUT116), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n690), .A2(KEYINPUT116), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n777), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n751), .A2(new_n685), .A3(new_n706), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n693), .A3(new_n715), .A4(new_n771), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n777), .A2(new_n778), .A3(new_n713), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n886), .A2(new_n770), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n886), .B2(new_n770), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n663), .A2(new_n427), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n891), .A2(new_n660), .A3(new_n662), .A4(new_n691), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n625), .A2(new_n783), .A3(new_n680), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n788), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n885), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n788), .A2(new_n893), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n797), .A2(new_n653), .A3(new_n714), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT114), .B1(new_n826), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n886), .A2(new_n770), .A3(new_n887), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n896), .A2(new_n900), .A3(KEYINPUT115), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n877), .A2(new_n884), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n693), .A2(new_n771), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n882), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n861), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT118), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n890), .A2(new_n885), .A3(new_n894), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT115), .B1(new_n896), .B2(new_n900), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n876), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n913));
  INV_X1    g727(.A(new_n907), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n884), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n906), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n740), .A2(new_n751), .A3(new_n493), .A4(new_n742), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n918), .A2(new_n831), .B1(new_n743), .B2(new_n666), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n749), .B1(new_n743), .B2(new_n650), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n902), .A2(new_n921), .A3(new_n872), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n882), .B(KEYINPUT52), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n907), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT119), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  INV_X1    g740(.A(new_n905), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n912), .A2(KEYINPUT53), .A3(new_n884), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n907), .C1(new_n922), .C2(new_n923), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n925), .A2(new_n926), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n917), .A2(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n860), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n707), .A2(new_n496), .A3(new_n364), .A4(new_n791), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n723), .B(KEYINPUT49), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n697), .A2(new_n935), .A3(new_n757), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n937), .ZN(G75));
  NOR2_X1   g752(.A1(new_n231), .A2(G952), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT122), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n925), .A2(new_n928), .A3(new_n930), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(G902), .ZN(new_n944));
  INV_X1    g758(.A(G210), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n535), .A2(new_n537), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n543), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT55), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n942), .B(new_n949), .C1(new_n944), .C2(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n951), .B2(new_n952), .ZN(G51));
  NAND2_X1  g767(.A1(new_n928), .A2(new_n930), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n929), .B1(new_n903), .B2(new_n907), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT54), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n931), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n355), .B(KEYINPUT123), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT57), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n352), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n944), .A2(new_n806), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n939), .B1(new_n960), .B2(new_n961), .ZN(G54));
  NAND2_X1  g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT124), .Z(new_n964));
  NAND3_X1  g778(.A1(new_n943), .A2(G902), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(new_n414), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n414), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n939), .ZN(G60));
  OR2_X1    g782(.A1(new_n644), .A2(new_n645), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT59), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n932), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n971), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n940), .B1(new_n957), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n954), .B2(new_n955), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n242), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(KEYINPUT125), .A3(new_n940), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n943), .A2(new_n678), .A3(new_n977), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n940), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n941), .B1(new_n978), .B2(new_n242), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n985), .B(new_n981), .C1(KEYINPUT125), .C2(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G66));
  INV_X1    g801(.A(G224), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n490), .B2(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n919), .A2(new_n920), .A3(new_n871), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n947), .B1(G898), .B2(new_n231), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  NAND4_X1  g807(.A1(new_n815), .A2(new_n699), .A3(new_n751), .A4(new_n852), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n904), .A2(new_n715), .ZN(new_n995));
  AND4_X1   g809(.A1(new_n786), .A2(new_n994), .A3(new_n788), .A4(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n816), .A2(new_n996), .A3(new_n231), .A4(new_n821), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n586), .B(new_n402), .Z(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n816), .A2(new_n821), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n995), .A2(new_n711), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n995), .A2(KEYINPUT62), .A3(new_n711), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n867), .A2(new_n700), .A3(new_n778), .ZN(new_n1006));
  AOI22_X1  g820(.A1(new_n1004), .A2(new_n1005), .B1(new_n734), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n998), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1000), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n231), .B1(G227), .B2(G900), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1011), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1000), .B(new_n1013), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(G72));
  NAND4_X1  g829(.A1(new_n816), .A2(new_n996), .A3(new_n821), .A4(new_n990), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n587), .B(KEYINPUT126), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1020), .A2(new_n578), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT127), .Z(new_n1022));
  AOI21_X1  g836(.A(new_n939), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n580), .A2(new_n616), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n916), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n816), .A2(new_n1007), .A3(new_n821), .A4(new_n990), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n1018), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1027), .A2(new_n578), .A3(new_n1020), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(G57));
endmodule


