

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573;

  XNOR2_X1 U317 ( .A(n398), .B(n397), .ZN(n515) );
  AND2_X1 U318 ( .A1(G230GAT), .A2(G233GAT), .ZN(n285) );
  XNOR2_X1 U319 ( .A(n360), .B(n285), .ZN(n342) );
  XNOR2_X1 U320 ( .A(n342), .B(n377), .ZN(n343) );
  XNOR2_X1 U321 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U322 ( .A(n396), .B(KEYINPUT48), .ZN(n397) );
  NOR2_X1 U323 ( .A1(n430), .A2(n514), .ZN(n431) );
  XNOR2_X1 U324 ( .A(n349), .B(n348), .ZN(n353) );
  NOR2_X1 U325 ( .A1(n447), .A2(n433), .ZN(n549) );
  XOR2_X1 U326 ( .A(n429), .B(n428), .Z(n514) );
  XNOR2_X1 U327 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n434) );
  XNOR2_X1 U328 ( .A(n435), .B(n434), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n287) );
  XNOR2_X1 U330 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n286) );
  XNOR2_X1 U331 ( .A(n287), .B(n286), .ZN(n288) );
  XOR2_X1 U332 ( .A(n288), .B(G183GAT), .Z(n290) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(G176GAT), .ZN(n289) );
  XNOR2_X1 U334 ( .A(n290), .B(n289), .ZN(n406) );
  XOR2_X1 U335 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n292) );
  NAND2_X1 U336 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n294) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G71GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n293), .B(G120GAT), .ZN(n351) );
  XOR2_X1 U340 ( .A(n294), .B(n351), .Z(n298) );
  XOR2_X1 U341 ( .A(G127GAT), .B(KEYINPUT82), .Z(n296) );
  XNOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n419) );
  XNOR2_X1 U344 ( .A(G15GAT), .B(n419), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n299), .B(KEYINPUT66), .Z(n301) );
  XOR2_X1 U347 ( .A(G43GAT), .B(G134GAT), .Z(n361) );
  XNOR2_X1 U348 ( .A(n361), .B(KEYINPUT83), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X2 U350 ( .A(n406), .B(n302), .Z(n517) );
  INV_X1 U351 ( .A(n517), .ZN(n447) );
  XOR2_X1 U352 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n304) );
  NAND2_X1 U353 ( .A1(G228GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U355 ( .A(n305), .B(KEYINPUT86), .Z(n310) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(KEYINPUT78), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n306), .B(G162GAT), .ZN(n364) );
  XOR2_X1 U358 ( .A(G155GAT), .B(KEYINPUT2), .Z(n308) );
  XNOR2_X1 U359 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n418) );
  XNOR2_X1 U361 ( .A(n364), .B(n418), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n316) );
  XOR2_X1 U363 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n314) );
  XOR2_X1 U364 ( .A(G78GAT), .B(G148GAT), .Z(n312) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n350) );
  XNOR2_X1 U367 ( .A(G204GAT), .B(n350), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n316), .B(n315), .Z(n322) );
  XNOR2_X1 U370 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n317), .B(KEYINPUT21), .ZN(n318) );
  XOR2_X1 U372 ( .A(n318), .B(KEYINPUT88), .Z(n320) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(G218GAT), .ZN(n319) );
  XOR2_X1 U374 ( .A(n320), .B(n319), .Z(n407) );
  XOR2_X1 U375 ( .A(G22GAT), .B(n407), .Z(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n448) );
  XOR2_X1 U377 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n411) );
  XOR2_X1 U378 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n355) );
  XOR2_X1 U379 ( .A(G113GAT), .B(G50GAT), .Z(n324) );
  XNOR2_X1 U380 ( .A(G169GAT), .B(G43GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U382 ( .A(KEYINPUT29), .B(n325), .Z(n327) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U385 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n329) );
  XNOR2_X1 U386 ( .A(G197GAT), .B(G141GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U388 ( .A(n331), .B(n330), .Z(n340) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n332), .B(G29GAT), .ZN(n333) );
  XOR2_X1 U391 ( .A(n333), .B(KEYINPUT71), .Z(n335) );
  XNOR2_X1 U392 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n359) );
  XOR2_X1 U394 ( .A(G22GAT), .B(G15GAT), .Z(n337) );
  XNOR2_X1 U395 ( .A(KEYINPUT72), .B(G1GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U397 ( .A(G8GAT), .B(n338), .Z(n376) );
  XNOR2_X1 U398 ( .A(n359), .B(n376), .ZN(n339) );
  XOR2_X1 U399 ( .A(n340), .B(n339), .Z(n490) );
  INV_X1 U400 ( .A(n490), .ZN(n554) );
  XOR2_X1 U401 ( .A(G92GAT), .B(G85GAT), .Z(n360) );
  XNOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n341), .B(KEYINPUT73), .ZN(n377) );
  XNOR2_X1 U404 ( .A(n343), .B(KEYINPUT74), .ZN(n349) );
  XOR2_X1 U405 ( .A(G204GAT), .B(G64GAT), .Z(n402) );
  XOR2_X1 U406 ( .A(G176GAT), .B(n402), .Z(n347) );
  XOR2_X1 U407 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n345) );
  XNOR2_X1 U408 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n344) );
  XOR2_X1 U409 ( .A(n345), .B(n344), .Z(n346) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n559) );
  XNOR2_X1 U412 ( .A(n559), .B(KEYINPUT41), .ZN(n542) );
  NAND2_X1 U413 ( .A1(n554), .A2(n542), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n389) );
  XOR2_X1 U415 ( .A(KEYINPUT9), .B(KEYINPUT67), .Z(n357) );
  XNOR2_X1 U416 ( .A(G99GAT), .B(KEYINPUT11), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n372) );
  XOR2_X1 U419 ( .A(KEYINPUT79), .B(n360), .Z(n363) );
  XNOR2_X1 U420 ( .A(n361), .B(G218GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U422 ( .A(n364), .B(KEYINPUT10), .Z(n366) );
  NAND2_X1 U423 ( .A1(G232GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U425 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U426 ( .A(G190GAT), .B(G106GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U428 ( .A(n372), .B(n371), .Z(n437) );
  INV_X1 U429 ( .A(n437), .ZN(n538) );
  XOR2_X1 U430 ( .A(KEYINPUT12), .B(G64GAT), .Z(n374) );
  XNOR2_X1 U431 ( .A(G155GAT), .B(G78GAT), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n387) );
  XOR2_X1 U434 ( .A(n377), .B(G211GAT), .Z(n379) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G71GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U437 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n381) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U440 ( .A(n383), .B(n382), .Z(n385) );
  XNOR2_X1 U441 ( .A(G183GAT), .B(KEYINPUT15), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U443 ( .A(n387), .B(n386), .Z(n472) );
  INV_X1 U444 ( .A(n472), .ZN(n563) );
  NOR2_X1 U445 ( .A1(n538), .A2(n563), .ZN(n388) );
  NAND2_X1 U446 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n390), .B(KEYINPUT47), .ZN(n395) );
  XOR2_X1 U448 ( .A(KEYINPUT36), .B(n538), .Z(n571) );
  NOR2_X1 U449 ( .A1(n571), .A2(n472), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT45), .ZN(n392) );
  NAND2_X1 U451 ( .A1(n392), .A2(n559), .ZN(n393) );
  NOR2_X1 U452 ( .A1(n393), .A2(n554), .ZN(n394) );
  NOR2_X1 U453 ( .A1(n395), .A2(n394), .ZN(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT64), .B(KEYINPUT112), .Z(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT92), .B(G92GAT), .Z(n400) );
  XNOR2_X1 U456 ( .A(G36GAT), .B(G8GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U458 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n409) );
  INV_X1 U462 ( .A(n407), .ZN(n408) );
  XOR2_X1 U463 ( .A(n409), .B(n408), .Z(n506) );
  NAND2_X1 U464 ( .A1(n515), .A2(n506), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n430) );
  XOR2_X1 U466 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n413) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(G57GAT), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n429) );
  XOR2_X1 U469 ( .A(G148GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U470 ( .A(G120GAT), .B(G134GAT), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U472 ( .A(G29GAT), .B(G85GAT), .Z(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n425) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n421) );
  XNOR2_X1 U476 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n427) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n431), .B(KEYINPUT65), .ZN(n553) );
  NOR2_X1 U483 ( .A1(n448), .A2(n553), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n432), .B(KEYINPUT55), .ZN(n433) );
  NAND2_X1 U485 ( .A1(n549), .A2(n538), .ZN(n435) );
  XOR2_X1 U486 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n460) );
  NAND2_X1 U487 ( .A1(n559), .A2(n554), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT77), .ZN(n476) );
  XOR2_X1 U489 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n439) );
  NAND2_X1 U490 ( .A1(n563), .A2(n437), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n458) );
  XNOR2_X1 U492 ( .A(n448), .B(KEYINPUT68), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n440), .B(KEYINPUT28), .ZN(n510) );
  XNOR2_X1 U494 ( .A(KEYINPUT27), .B(KEYINPUT93), .ZN(n441) );
  INV_X1 U495 ( .A(n506), .ZN(n444) );
  XOR2_X1 U496 ( .A(n441), .B(n444), .Z(n452) );
  NOR2_X1 U497 ( .A1(n510), .A2(n452), .ZN(n516) );
  XNOR2_X1 U498 ( .A(KEYINPUT85), .B(n517), .ZN(n442) );
  NAND2_X1 U499 ( .A1(n516), .A2(n442), .ZN(n443) );
  NAND2_X1 U500 ( .A1(n443), .A2(n514), .ZN(n457) );
  NOR2_X1 U501 ( .A1(n444), .A2(n447), .ZN(n445) );
  NOR2_X1 U502 ( .A1(n448), .A2(n445), .ZN(n446) );
  XNOR2_X1 U503 ( .A(KEYINPUT25), .B(n446), .ZN(n455) );
  XOR2_X1 U504 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n450) );
  NAND2_X1 U505 ( .A1(n448), .A2(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT94), .B(n451), .ZN(n552) );
  OR2_X1 U508 ( .A1(n552), .A2(n452), .ZN(n530) );
  XOR2_X1 U509 ( .A(KEYINPUT96), .B(n530), .Z(n453) );
  NOR2_X1 U510 ( .A1(n514), .A2(n453), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n457), .A2(n456), .ZN(n471) );
  NOR2_X1 U513 ( .A1(n458), .A2(n471), .ZN(n491) );
  AND2_X1 U514 ( .A1(n476), .A2(n491), .ZN(n467) );
  NAND2_X1 U515 ( .A1(n467), .A2(n514), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U517 ( .A(G1GAT), .B(n461), .ZN(G1324GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n463) );
  NAND2_X1 U519 ( .A1(n467), .A2(n506), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U521 ( .A(G8GAT), .B(n464), .ZN(G1325GAT) );
  XOR2_X1 U522 ( .A(G15GAT), .B(KEYINPUT35), .Z(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n517), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(G1326GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n469) );
  NAND2_X1 U526 ( .A1(n467), .A2(n510), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(G22GAT), .B(n470), .ZN(G1327GAT) );
  XNOR2_X1 U529 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n571), .A2(n471), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U532 ( .A(n475), .B(n474), .Z(n504) );
  INV_X1 U533 ( .A(n504), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n480) );
  XNOR2_X1 U535 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT104), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n487), .A2(n514), .ZN(n483) );
  XNOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT39), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1328GAT) );
  NAND2_X1 U542 ( .A1(n506), .A2(n487), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U544 ( .A1(n517), .A2(n487), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT40), .B(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(G43GAT), .B(n486), .ZN(G1330GAT) );
  NAND2_X1 U547 ( .A1(n487), .A2(n510), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT106), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G50GAT), .B(n489), .ZN(G1331GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n494) );
  NAND2_X1 U551 ( .A1(n490), .A2(n542), .ZN(n503) );
  INV_X1 U552 ( .A(n491), .ZN(n492) );
  NOR2_X1 U553 ( .A1(n503), .A2(n492), .ZN(n499) );
  NAND2_X1 U554 ( .A1(n499), .A2(n514), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(n495), .ZN(G1332GAT) );
  NAND2_X1 U557 ( .A1(n506), .A2(n499), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U559 ( .A1(n499), .A2(n517), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT108), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G71GAT), .B(n498), .ZN(G1334GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n501) );
  NAND2_X1 U563 ( .A1(n499), .A2(n510), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U565 ( .A(G78GAT), .B(n502), .Z(G1335GAT) );
  NOR2_X1 U566 ( .A1(n504), .A2(n503), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n511), .A2(n514), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U569 ( .A1(n506), .A2(n511), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U571 ( .A1(n511), .A2(n517), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G99GAT), .B(n509), .ZN(G1338GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(KEYINPUT44), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G106GAT), .B(n513), .ZN(G1339GAT) );
  XOR2_X1 U577 ( .A(G113GAT), .B(KEYINPUT113), .Z(n520) );
  NAND2_X1 U578 ( .A1(n515), .A2(n514), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U580 ( .A1(n529), .A2(n518), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n526), .A2(n554), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1340GAT) );
  XOR2_X1 U583 ( .A(G120GAT), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U584 ( .A1(n526), .A2(n542), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1341GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n524) );
  NAND2_X1 U587 ( .A1(n526), .A2(n563), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U589 ( .A(G127GAT), .B(n525), .Z(G1342GAT) );
  XOR2_X1 U590 ( .A(G134GAT), .B(KEYINPUT51), .Z(n528) );
  NAND2_X1 U591 ( .A1(n526), .A2(n538), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1343GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n554), .A2(n539), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G141GAT), .B(n531), .ZN(G1344GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT53), .Z(n533) );
  NAND2_X1 U597 ( .A1(n539), .A2(n542), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U599 ( .A(G148GAT), .B(KEYINPUT52), .Z(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1345GAT) );
  NAND2_X1 U601 ( .A1(n539), .A2(n563), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT116), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G155GAT), .B(n537), .ZN(G1346GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U606 ( .A1(n554), .A2(n549), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G169GAT), .B(n541), .ZN(G1348GAT) );
  NAND2_X1 U608 ( .A1(n542), .A2(n549), .ZN(n548) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n544) );
  XNOR2_X1 U610 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U612 ( .A(G176GAT), .B(KEYINPUT118), .Z(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1349GAT) );
  XOR2_X1 U615 ( .A(G183GAT), .B(KEYINPUT121), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n563), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1350GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n564), .A2(n554), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n556) );
  XNOR2_X1 U621 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1352GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n561) );
  INV_X1 U625 ( .A(n564), .ZN(n570) );
  OR2_X1 U626 ( .A1(n570), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G204GAT), .B(n562), .Z(G1353GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n566) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G211GAT), .B(n567), .ZN(G1354GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n569) );
  XNOR2_X1 U634 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(n573), .B(n572), .Z(G1355GAT) );
endmodule

