//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1182, new_n1183,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AND2_X1   g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G87), .C2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G50), .A2(G226), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n209), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT64), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT7), .ZN(new_n250));
  NOR3_X1   g0050(.A1(new_n249), .A2(new_n250), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT7), .B1(new_n256), .B2(new_n227), .ZN(new_n257));
  OAI21_X1  g0057(.A(G68), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n227), .A2(new_n252), .A3(G159), .ZN(new_n259));
  INV_X1    g0059(.A(G58), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n221), .ZN(new_n261));
  OAI21_X1  g0061(.A(G20), .B1(new_n261), .B2(new_n201), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT16), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n226), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n258), .A2(KEYINPUT16), .A3(new_n259), .A4(new_n262), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT8), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(new_n271), .A3(G58), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT68), .B1(new_n271), .B2(G58), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n260), .A2(KEYINPUT8), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n277), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n267), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G1), .B2(new_n227), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n276), .A3(new_n278), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n269), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT66), .A2(G41), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT66), .A2(G41), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n280), .B(G274), .C1(new_n292), .C2(G45), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n280), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n252), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n280), .C1(G41), .C2(G45), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G232), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n293), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(G226), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n249), .B(new_n304), .C1(G223), .C2(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G87), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n297), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n289), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n302), .A2(new_n307), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT70), .B(G179), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n288), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT18), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n288), .A2(KEYINPUT18), .A3(new_n308), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n309), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(G200), .B2(new_n309), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n319), .A2(new_n269), .A3(new_n283), .A4(new_n287), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT74), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n320), .B1(new_n323), .B2(KEYINPUT17), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n281), .A2(G77), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G20), .A2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n227), .A2(G33), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n227), .A2(new_n252), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n327), .B1(new_n328), .B2(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(new_n332), .B2(new_n267), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n211), .B2(new_n285), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT71), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n249), .A2(G232), .A3(new_n303), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n256), .A2(G107), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n297), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n300), .A2(new_n212), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(new_n293), .A3(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n334), .B(new_n335), .C1(new_n343), .C2(G169), .ZN(new_n344));
  INV_X1    g0144(.A(new_n293), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n339), .B2(new_n340), .ZN(new_n346));
  AOI21_X1  g0146(.A(G169), .B1(new_n346), .B2(new_n342), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n211), .B(new_n267), .C1(new_n280), .C2(G20), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n326), .B(new_n348), .C1(new_n267), .C2(new_n332), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT71), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n343), .A2(new_n310), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(G190), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n349), .C1(new_n354), .C2(new_n343), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n316), .A2(new_n325), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n293), .B1(new_n300), .B2(new_n222), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n301), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n249), .B(new_n359), .C1(G226), .C2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n297), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR3_X1    g0162(.A1(new_n358), .A2(new_n362), .A3(KEYINPUT13), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT13), .B1(new_n358), .B2(new_n362), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n289), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(G179), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n366), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n331), .A2(new_n202), .B1(new_n227), .B2(G68), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n329), .A2(new_n211), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n267), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g0173(.A(new_n373), .B(KEYINPUT11), .Z(new_n374));
  INV_X1    g0174(.A(KEYINPUT12), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n282), .B2(new_n221), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n285), .A2(new_n221), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n363), .A2(new_n364), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(G200), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n317), .B2(new_n382), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n203), .A2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n227), .A2(new_n252), .A3(G150), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n386), .B(new_n387), .C1(new_n279), .C2(new_n329), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n267), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n285), .A2(new_n202), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n281), .A2(G50), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(G222), .A2(G1698), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n303), .A2(G223), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n249), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n340), .C1(G77), .C2(new_n249), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n295), .A2(G226), .A3(new_n297), .A4(new_n299), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n293), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n289), .ZN(new_n401));
  INV_X1    g0201(.A(new_n310), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n394), .B(new_n401), .C1(new_n402), .C2(new_n400), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n398), .A2(G190), .A3(new_n293), .A4(new_n399), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT73), .ZN(new_n405));
  AOI211_X1 g0205(.A(new_n390), .B(new_n392), .C1(new_n388), .C2(new_n267), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(KEYINPUT9), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(G200), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT72), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n406), .A2(new_n409), .A3(KEYINPUT9), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT9), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT72), .B1(new_n394), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n407), .B(new_n408), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n409), .B1(new_n406), .B2(KEYINPUT9), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n394), .A2(KEYINPUT72), .A3(new_n411), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT10), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n408), .A4(new_n407), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  AND4_X1   g0220(.A1(new_n357), .A2(new_n385), .A3(new_n403), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G116), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n282), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n280), .A2(G33), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n284), .A2(G116), .A3(new_n281), .A4(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n266), .A2(new_n226), .B1(G20), .B2(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G283), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n227), .C1(G33), .C2(new_n213), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n426), .A2(KEYINPUT20), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT20), .B1(new_n426), .B2(new_n428), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n423), .B(new_n425), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n254), .A2(G33), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n434));
  OAI21_X1  g0234(.A(G303), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n253), .A2(new_n255), .A3(G257), .A4(new_n303), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n253), .A2(new_n255), .A3(G264), .A4(G1698), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n340), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT5), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT5), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n280), .B(G45), .C1(new_n441), .C2(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n297), .B(G270), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n442), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT66), .A2(G41), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT66), .A2(G41), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n444), .B(G274), .C1(KEYINPUT5), .C2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n439), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT21), .A3(G169), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n439), .A2(G179), .A3(new_n443), .A4(new_n448), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n432), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n438), .A2(new_n340), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n443), .A2(new_n448), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n431), .B(G169), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT21), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(KEYINPUT77), .A3(new_n456), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n452), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(new_n303), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n249), .A2(KEYINPUT80), .A3(G250), .A4(new_n303), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n253), .A2(new_n255), .A3(G257), .A4(G1698), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G294), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT81), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT81), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(new_n464), .A4(new_n465), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n340), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n297), .B(G264), .C1(new_n440), .C2(new_n442), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n448), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n289), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT23), .B1(new_n227), .B2(G107), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  INV_X1    g0280(.A(G107), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(G20), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n479), .A2(new_n482), .A3(new_n483), .A4(KEYINPUT79), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n253), .A2(new_n255), .A3(new_n227), .A4(G87), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT22), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n489), .B(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n478), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n486), .A2(new_n487), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n490), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n489), .A2(new_n490), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(KEYINPUT24), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n267), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n281), .A2(new_n424), .A3(new_n226), .A4(new_n266), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G107), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n281), .A2(G107), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT25), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G179), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n474), .A2(new_n504), .A3(new_n475), .A4(new_n448), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n477), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n461), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n253), .A2(new_n255), .A3(G244), .A4(new_n303), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n303), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n427), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n340), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n297), .B(G257), .C1(new_n440), .C2(new_n442), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n516), .A2(new_n448), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n517), .A3(new_n310), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT76), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n517), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n289), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n522), .A2(new_n213), .A3(G107), .ZN(new_n523));
  XNOR2_X1  g0323(.A(G97), .B(G107), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n525), .A2(new_n227), .B1(new_n211), .B2(new_n331), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n250), .B1(new_n249), .B2(G20), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n481), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n267), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n499), .A2(G97), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n282), .A2(new_n213), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n532), .B(KEYINPUT75), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT76), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n515), .A2(new_n517), .A3(new_n535), .A4(new_n310), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n519), .A2(new_n521), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n520), .A2(G200), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n331), .A2(new_n211), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n524), .A2(new_n522), .ZN(new_n540));
  INV_X1    g0340(.A(new_n523), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n542), .B2(G20), .ZN(new_n543));
  OAI21_X1  g0343(.A(G107), .B1(new_n251), .B2(new_n257), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n267), .B1(G97), .B2(new_n499), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n515), .A2(new_n517), .A3(G190), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n538), .A2(new_n546), .A3(new_n533), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n227), .ZN(new_n550));
  INV_X1    g0350(.A(G87), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n213), .A3(new_n481), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n227), .A2(G33), .A3(G97), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n550), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n253), .A2(new_n255), .A3(new_n227), .A4(G68), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n284), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n328), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n281), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n498), .A2(new_n551), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n222), .A2(new_n303), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n212), .A2(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n253), .A2(new_n562), .A3(new_n255), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n340), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n280), .A2(G45), .A3(G274), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n280), .A2(G45), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n297), .A2(G250), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n567), .A2(G190), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n297), .B1(new_n564), .B2(new_n565), .ZN(new_n572));
  INV_X1    g0372(.A(new_n570), .ZN(new_n573));
  INV_X1    g0373(.A(new_n568), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n561), .B(new_n571), .C1(new_n575), .C2(new_n354), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n550), .A2(new_n552), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n553), .A2(new_n554), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n556), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n267), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n499), .A2(new_n558), .ZN(new_n581));
  INV_X1    g0381(.A(new_n559), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n567), .A2(new_n310), .A3(new_n568), .A4(new_n570), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n575), .C2(G169), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n537), .A2(new_n548), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n474), .A2(G190), .A3(new_n475), .A4(new_n448), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n503), .B1(G200), .B2(new_n476), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n453), .A2(new_n454), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n432), .B1(new_n591), .B2(new_n354), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT78), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n421), .A2(new_n508), .A3(new_n590), .A4(new_n597), .ZN(G372));
  INV_X1    g0398(.A(new_n403), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n414), .A2(KEYINPUT84), .A3(new_n419), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT84), .B1(new_n414), .B2(new_n419), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n352), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n344), .A2(new_n350), .A3(KEYINPUT83), .A4(new_n351), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n384), .B1(new_n370), .B2(new_n380), .ZN(new_n607));
  INV_X1    g0407(.A(new_n325), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n316), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n599), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n385), .A2(new_n420), .A3(new_n403), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n357), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n476), .A2(G200), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n613), .A2(new_n588), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT82), .B1(new_n615), .B2(new_n587), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n537), .A2(new_n548), .A3(new_n586), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT82), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n588), .A3(new_n614), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n616), .A2(new_n507), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n585), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n519), .A2(new_n536), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n521), .A2(new_n534), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n586), .A4(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n576), .A2(new_n585), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n537), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n610), .B1(new_n612), .B2(new_n630), .ZN(G369));
  INV_X1    g0431(.A(new_n461), .ZN(new_n632));
  INV_X1    g0432(.A(new_n597), .ZN(new_n633));
  INV_X1    g0433(.A(G13), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n280), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(KEYINPUT85), .B(G343), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT86), .Z(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n432), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n632), .B1(new_n633), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT87), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n619), .B1(new_n613), .B2(new_n642), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n506), .ZN(new_n653));
  INV_X1    g0453(.A(new_n642), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n506), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n461), .A2(new_n654), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n207), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n292), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n552), .A2(G116), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G1), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n229), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n507), .A2(new_n617), .A3(new_n619), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n629), .ZN(new_n669));
  AND4_X1   g0469(.A1(KEYINPUT89), .A2(new_n669), .A3(KEYINPUT29), .A4(new_n642), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n654), .B1(new_n668), .B2(new_n629), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT89), .B1(new_n671), .B2(KEYINPUT29), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n654), .B1(new_n621), .B2(new_n629), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n670), .A2(new_n672), .B1(new_n673), .B2(KEYINPUT29), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n590), .A2(new_n508), .A3(new_n597), .A4(new_n642), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n474), .A2(new_n475), .ZN(new_n676));
  INV_X1    g0476(.A(new_n451), .ZN(new_n677));
  INV_X1    g0477(.A(new_n575), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n520), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n676), .A2(KEYINPUT30), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n516), .A2(new_n448), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n340), .B2(new_n514), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n474), .A2(new_n683), .A3(new_n475), .A4(new_n575), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n681), .B1(new_n684), .B2(new_n451), .ZN(new_n685));
  INV_X1    g0485(.A(new_n476), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n678), .A2(KEYINPUT88), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT88), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n402), .B1(new_n575), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n687), .A2(new_n689), .A3(new_n449), .A4(new_n520), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n680), .B(new_n685), .C1(new_n686), .C2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n654), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n675), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n674), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n667), .B1(new_n699), .B2(G1), .ZN(G364));
  NAND2_X1  g0500(.A1(new_n635), .A2(G45), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n663), .A2(G1), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n651), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(G330), .B2(new_n650), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n661), .A2(new_n249), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n243), .B2(G45), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(G45), .B2(new_n229), .ZN(new_n709));
  INV_X1    g0509(.A(G355), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n249), .A2(new_n207), .ZN(new_n711));
  OAI221_X1 g0511(.A(new_n709), .B1(G116), .B2(new_n207), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n226), .B1(G20), .B2(new_n289), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n227), .A2(G179), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G190), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G159), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT32), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n310), .A2(new_n227), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n317), .A2(new_n354), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n249), .B1(new_n730), .B2(new_n202), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n317), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n724), .B(new_n731), .C1(G58), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n354), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G107), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n725), .A2(new_n720), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G77), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n227), .B1(new_n732), .B2(new_n504), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n213), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n727), .A2(new_n719), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n551), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n725), .A2(new_n736), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n744), .B(new_n746), .C1(new_n748), .C2(G68), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n735), .A2(new_n739), .A3(new_n742), .A4(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G322), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n733), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n743), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n729), .A2(G326), .B1(G294), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n755), .A2(KEYINPUT90), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G283), .A2(new_n738), .B1(new_n722), .B2(G329), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n256), .C1(new_n759), .C2(new_n745), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT90), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(new_n754), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n757), .B(new_n762), .C1(new_n763), .C2(new_n740), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n750), .B1(new_n752), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n716), .ZN(new_n766));
  INV_X1    g0566(.A(new_n715), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n718), .B(new_n766), .C1(new_n650), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n705), .B1(new_n702), .B2(new_n768), .ZN(G396));
  NAND2_X1  g0569(.A1(new_n654), .A2(new_n334), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n356), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n604), .A2(new_n605), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n772), .B2(new_n770), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n673), .B(new_n773), .Z(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(new_n697), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n702), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n730), .A2(new_n759), .B1(new_n422), .B2(new_n740), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G283), .B2(new_n748), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT92), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n745), .A2(new_n481), .B1(new_n737), .B2(new_n551), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n779), .A2(new_n249), .A3(new_n744), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n781), .B1(new_n782), .B2(new_n733), .C1(new_n763), .C2(new_n721), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n745), .A2(new_n202), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n737), .A2(new_n221), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G143), .A2(new_n734), .B1(new_n741), .B2(G159), .ZN(new_n787));
  INV_X1    g0587(.A(G137), .ZN(new_n788));
  INV_X1    g0588(.A(G150), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n788), .B2(new_n730), .C1(new_n789), .C2(new_n747), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n785), .B(new_n786), .C1(new_n791), .C2(KEYINPUT34), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n753), .A2(G58), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n256), .B1(new_n722), .B2(G132), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT34), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n790), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n716), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n716), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n714), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n211), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n773), .A2(new_n714), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n798), .A2(new_n703), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n776), .A2(new_n804), .ZN(G384));
  INV_X1    g0605(.A(KEYINPUT38), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n288), .A2(new_n639), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n312), .A2(new_n320), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT37), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT37), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n312), .A2(new_n807), .A3(new_n810), .A4(new_n320), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n807), .B1(new_n316), .B2(new_n325), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n809), .A2(new_n811), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n316), .A2(new_n325), .ZN(new_n816));
  OAI211_X1 g0616(.A(KEYINPUT38), .B(new_n815), .C1(new_n816), .C2(new_n807), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n642), .A2(new_n379), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n370), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n381), .A2(new_n384), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n819), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n696), .A2(new_n822), .A3(new_n773), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT40), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G330), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n611), .A2(new_n696), .A3(new_n357), .A4(G330), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT96), .Z(new_n829));
  NAND3_X1  g0629(.A1(new_n825), .A2(new_n421), .A3(new_n696), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n673), .A2(KEYINPUT29), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT89), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n671), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n832), .A2(new_n837), .A3(new_n421), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n610), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n831), .B(new_n839), .Z(new_n840));
  NOR2_X1   g0640(.A1(new_n316), .A2(new_n639), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT94), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT95), .Z(new_n844));
  NOR2_X1   g0644(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n818), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n844), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n845), .B(new_n848), .C1(new_n814), .C2(new_n817), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n381), .A2(new_n654), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n841), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n352), .A2(new_n654), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n673), .B2(new_n773), .ZN(new_n854));
  INV_X1    g0654(.A(new_n822), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n818), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n840), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n280), .B2(new_n635), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n422), .B1(new_n542), .B2(KEYINPUT35), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n861), .B(new_n228), .C1(KEYINPUT35), .C2(new_n542), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT36), .ZN(new_n863));
  OAI21_X1  g0663(.A(G77), .B1(new_n260), .B2(new_n221), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n864), .A2(new_n229), .B1(G50), .B2(new_n221), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(G1), .A3(new_n634), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n860), .A2(new_n863), .A3(new_n866), .ZN(G367));
  OAI22_X1  g0667(.A1(new_n730), .A2(new_n763), .B1(new_n782), .B2(new_n747), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n249), .B(new_n868), .C1(G303), .C2(new_n734), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n745), .A2(new_n422), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n870), .A2(KEYINPUT46), .B1(new_n481), .B2(new_n743), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(KEYINPUT46), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n213), .B2(new_n737), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n871), .B(new_n873), .C1(G317), .C2(new_n722), .ZN(new_n874));
  INV_X1    g0674(.A(G283), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n869), .B(new_n874), .C1(new_n875), .C2(new_n740), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n202), .A2(new_n740), .B1(new_n733), .B2(new_n789), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G143), .B2(new_n729), .ZN(new_n878));
  INV_X1    g0678(.A(G159), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n747), .A2(new_n879), .B1(new_n221), .B2(new_n743), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n249), .B1(new_n737), .B2(new_n211), .C1(new_n260), .C2(new_n745), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n878), .B(new_n882), .C1(new_n788), .C2(new_n721), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT47), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n716), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n642), .A2(new_n561), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(new_n586), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n715), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n717), .B1(new_n207), .B2(new_n328), .C1(new_n238), .C2(new_n707), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n886), .A2(new_n703), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n701), .A2(G1), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n650), .A2(G330), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n656), .A2(new_n658), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n656), .A2(new_n658), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(KEYINPUT103), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n699), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n654), .A2(new_n534), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n537), .A2(new_n548), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n642), .A2(new_n537), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n659), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT45), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT100), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n659), .A2(KEYINPUT45), .A3(new_n906), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n901), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n909), .A2(new_n911), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(KEYINPUT101), .A3(new_n912), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n659), .A2(new_n906), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT44), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n915), .A2(new_n918), .A3(new_n657), .A4(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n921), .A2(new_n922), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n900), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n915), .A2(new_n918), .A3(new_n920), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT102), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n657), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT102), .A4(new_n920), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n926), .A2(new_n933), .A3(KEYINPUT105), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n921), .A2(new_n922), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n899), .B1(new_n936), .B2(new_n923), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n935), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n699), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n662), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n892), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n896), .A2(new_n903), .A3(new_n902), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT97), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n537), .B1(new_n904), .B2(new_n506), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n642), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT98), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n888), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n888), .A2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n954), .A3(new_n888), .A4(new_n952), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n930), .A2(new_n906), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n891), .B1(new_n943), .B2(new_n961), .ZN(G387));
  AOI22_X1  g0762(.A1(G322), .A2(new_n729), .B1(new_n748), .B2(G311), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n759), .B2(new_n740), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G317), .B2(new_n734), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT48), .Z(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n875), .B2(new_n743), .C1(new_n782), .C2(new_n745), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT108), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT49), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n249), .B1(new_n722), .B2(G326), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n970), .C1(new_n422), .C2(new_n737), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n249), .B1(new_n279), .B2(new_n747), .C1(new_n730), .C2(new_n879), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G50), .B2(new_n734), .ZN(new_n973));
  INV_X1    g0773(.A(new_n745), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(G77), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n741), .A2(G68), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n743), .A2(new_n328), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n789), .B2(new_n721), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G97), .B2(new_n738), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n973), .A2(new_n975), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n799), .B1(new_n971), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n330), .A2(G50), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT50), .ZN(new_n984));
  AOI211_X1 g0784(.A(G116), .B(new_n552), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(G45), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n984), .C2(new_n983), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n221), .A2(new_n211), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n706), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n986), .B2(new_n235), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n711), .A2(new_n664), .B1(G107), .B2(new_n207), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT106), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n702), .B(new_n982), .C1(new_n717), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n656), .B2(new_n767), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n898), .A2(new_n892), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n662), .B1(new_n898), .B2(new_n699), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n997), .C1(new_n900), .C2(new_n998), .ZN(G393));
  AOI22_X1  g0799(.A1(G68), .A2(new_n974), .B1(new_n722), .B2(G143), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n1000), .A2(KEYINPUT109), .B1(new_n202), .B2(new_n747), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n730), .A2(new_n789), .B1(new_n879), .B2(new_n733), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT51), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n743), .A2(new_n211), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n256), .B(new_n1004), .C1(G87), .C2(new_n738), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(new_n330), .C2(new_n740), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1001), .B(new_n1006), .C1(KEYINPUT109), .C2(new_n1000), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G317), .A2(new_n729), .B1(new_n734), .B2(G311), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1008), .A2(new_n1010), .B1(new_n759), .B2(new_n747), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n739), .B1(new_n751), .B2(new_n721), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n249), .B(new_n1012), .C1(G116), .C2(new_n753), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n782), .C2(new_n740), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1011), .B(new_n1015), .C1(G283), .C2(new_n974), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n716), .B1(new_n1007), .B2(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n717), .B1(new_n213), .B2(new_n207), .C1(new_n247), .C2(new_n707), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n904), .A2(new_n715), .A3(new_n905), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1017), .A2(new_n703), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n927), .A2(new_n930), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n924), .B2(new_n925), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n892), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT105), .B1(new_n926), .B2(new_n933), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n937), .A2(new_n935), .A3(new_n932), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1025), .A2(new_n1026), .B1(new_n899), .B2(new_n1022), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1027), .B2(new_n662), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G390));
  OAI22_X1  g0829(.A1(new_n847), .A2(new_n849), .B1(new_n856), .B2(new_n851), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n696), .A2(new_n822), .A3(G330), .A4(new_n773), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT111), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n773), .A2(new_n671), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n853), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n822), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n851), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n818), .A3(new_n1039), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1030), .A2(new_n1031), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1031), .B1(new_n1030), .B2(new_n1040), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n696), .A2(G330), .A3(new_n773), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n855), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1031), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n854), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1037), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1045), .B(new_n1031), .C1(new_n1049), .C2(new_n1035), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n610), .B(new_n827), .C1(new_n674), .C2(new_n612), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n838), .A2(new_n1054), .A3(new_n610), .A4(new_n827), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT113), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT113), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1051), .A2(new_n1053), .A3(new_n1058), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT114), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1060), .A2(new_n1043), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1060), .B2(new_n1043), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n662), .B1(new_n1043), .B2(new_n1060), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1043), .A2(new_n892), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n713), .B1(new_n847), .B2(new_n849), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1004), .B1(new_n729), .B2(G283), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT117), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n213), .A2(new_n740), .B1(new_n747), .B2(new_n481), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n786), .B(new_n1070), .C1(G116), .C2(new_n734), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n256), .B1(new_n721), .B2(new_n782), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n746), .B(new_n1072), .C1(new_n1069), .C2(new_n1068), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G128), .ZN(new_n1075));
  INV_X1    g0875(.A(G132), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n730), .A2(new_n1075), .B1(new_n1076), .B2(new_n733), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT116), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n748), .A2(G137), .ZN(new_n1079));
  INV_X1    g0879(.A(G125), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n743), .A2(new_n879), .B1(new_n721), .B2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT115), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n256), .B(new_n1081), .C1(new_n741), .C2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n974), .A2(G150), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(KEYINPUT53), .B1(new_n738), .B2(G50), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1078), .A2(new_n1079), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1085), .A2(KEYINPUT53), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1074), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n716), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n801), .A2(new_n279), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1066), .A2(new_n703), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1064), .A2(new_n1065), .A3(new_n1092), .ZN(G378));
  INV_X1    g0893(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1060), .A2(new_n1043), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT114), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1060), .A2(new_n1043), .A3(new_n1061), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n394), .A2(new_n639), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n602), .B2(new_n403), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1103));
  NAND3_X1  g0903(.A1(new_n602), .A2(new_n403), .A3(new_n1100), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n826), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n826), .A2(new_n1107), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n858), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n857), .A3(new_n852), .A4(new_n1109), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1094), .B1(new_n1099), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1095), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1112), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1108), .A2(new_n1109), .B1(new_n852), .B2(new_n857), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1119), .A3(KEYINPUT57), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1114), .A2(new_n662), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n892), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n713), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n730), .A2(new_n422), .B1(new_n213), .B2(new_n747), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n558), .B2(new_n741), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n975), .A2(new_n256), .A3(new_n447), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n733), .A2(new_n481), .B1(new_n221), .B2(new_n743), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(G283), .C2(new_n722), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1129), .C1(new_n260), .C2(new_n737), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(G33), .A2(G41), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n202), .B1(new_n292), .B2(new_n249), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n734), .A2(G128), .B1(new_n1083), .B2(new_n974), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT119), .Z(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n1076), .B2(new_n747), .C1(new_n788), .C2(new_n740), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G150), .B2(new_n753), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1080), .B2(new_n730), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT59), .ZN(new_n1140));
  INV_X1    g0940(.A(G124), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1133), .B1(new_n721), .B2(new_n1141), .C1(new_n879), .C2(new_n737), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n716), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n801), .A2(new_n202), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1124), .A2(new_n703), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1123), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1121), .A2(new_n1122), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1122), .B1(new_n1121), .B2(new_n1147), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G375));
  NAND2_X1  g0952(.A1(new_n855), .A2(new_n713), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n801), .A2(new_n221), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n729), .A2(G132), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT122), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n249), .B1(new_n733), .B2(new_n788), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n740), .A2(new_n789), .B1(new_n1075), .B2(new_n721), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G58), .C2(new_n738), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n974), .A2(G159), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n748), .A2(new_n1083), .B1(G50), .B2(new_n753), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1157), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n747), .A2(new_n422), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n978), .B1(new_n733), .B2(new_n875), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT121), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n741), .A2(G107), .B1(G97), .B2(new_n974), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n737), .A2(new_n211), .B1(new_n721), .B2(new_n759), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n249), .B(new_n1168), .C1(new_n729), .C2(G294), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1163), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n702), .B(new_n1155), .C1(new_n716), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1051), .B2(new_n892), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1095), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1057), .A2(new_n1174), .A3(new_n1059), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1175), .B2(new_n941), .ZN(G381));
  INV_X1    g0976(.A(G378), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(G381), .A2(G384), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1151), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n891), .B(new_n1028), .C1(new_n943), .C2(new_n961), .ZN(new_n1180));
  OR4_X1    g0980(.A1(G396), .A2(new_n1179), .A3(G393), .A4(new_n1180), .ZN(G407));
  INV_X1    g0981(.A(new_n640), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1151), .A2(new_n1182), .A3(new_n1177), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(G407), .A2(G213), .A3(new_n1183), .ZN(G409));
  INV_X1    g0984(.A(KEYINPUT62), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT124), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1113), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1111), .A2(KEYINPUT124), .A3(new_n1112), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n892), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1116), .A2(new_n1119), .A3(new_n942), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1146), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1177), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1121), .A2(G378), .A3(new_n1147), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT123), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1121), .A2(G378), .A3(new_n1196), .A4(new_n1147), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1193), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1182), .A2(G213), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  MUX2_X1   g1000(.A(new_n1174), .B(new_n1175), .S(KEYINPUT60), .Z(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(new_n663), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1173), .ZN(new_n1203));
  INV_X1    g1003(.A(G384), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(G384), .A3(new_n1173), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1198), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT125), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1185), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1192), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1207), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1199), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1199), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1200), .A2(G2897), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1207), .B(new_n1217), .Z(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT61), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1210), .A2(new_n1215), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(G387), .A2(G390), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(G393), .B(G396), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1222), .A2(new_n1180), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1222), .B2(new_n1180), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1218), .B1(new_n1199), .B2(new_n1212), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT63), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1214), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1208), .A2(KEYINPUT63), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1226), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1228), .A2(new_n1234), .ZN(G405));
  OAI21_X1  g1035(.A(new_n1177), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1213), .A2(KEYINPUT126), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1211), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1237), .B1(new_n1236), .B2(new_n1211), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT127), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1211), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1213), .A2(KEYINPUT126), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1238), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1241), .A2(new_n1226), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1226), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(G402));
endmodule


