

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734;

  INV_X1 U357 ( .A(G953), .ZN(n726) );
  XNOR2_X2 U358 ( .A(n435), .B(n434), .ZN(n707) );
  NOR2_X2 U359 ( .A1(n601), .A2(n571), .ZN(n572) );
  NOR2_X2 U360 ( .A1(n548), .A2(n539), .ZN(n540) );
  XNOR2_X1 U361 ( .A(G104), .B(G110), .ZN(n475) );
  XNOR2_X1 U362 ( .A(G116), .B(G113), .ZN(n479) );
  NOR2_X2 U363 ( .A1(G953), .A2(G237), .ZN(n520) );
  NAND2_X1 U364 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U365 ( .A1(n442), .A2(n436), .ZN(n547) );
  AND2_X1 U366 ( .A1(n597), .A2(n363), .ZN(n362) );
  AND2_X1 U367 ( .A1(n593), .A2(n592), .ZN(n632) );
  XNOR2_X1 U368 ( .A(n583), .B(KEYINPUT39), .ZN(n611) );
  NOR2_X1 U369 ( .A1(n607), .A2(n603), .ZN(n604) );
  NAND2_X2 U370 ( .A1(n390), .A2(n388), .ZN(n558) );
  NAND2_X1 U371 ( .A1(n389), .A2(n338), .ZN(n388) );
  AND2_X1 U372 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U373 ( .A1(n503), .A2(n393), .ZN(n391) );
  XNOR2_X1 U374 ( .A(n471), .B(n470), .ZN(n702) );
  XNOR2_X1 U375 ( .A(n474), .B(KEYINPUT25), .ZN(n430) );
  XNOR2_X1 U376 ( .A(n479), .B(n481), .ZN(n449) );
  XNOR2_X1 U377 ( .A(n475), .B(G107), .ZN(n532) );
  NAND2_X1 U378 ( .A1(n365), .A2(n389), .ZN(n633) );
  NOR2_X1 U379 ( .A1(n732), .A2(n627), .ZN(n541) );
  XNOR2_X1 U380 ( .A(n379), .B(n525), .ZN(n415) );
  XNOR2_X2 U381 ( .A(n431), .B(n519), .ZN(n710) );
  XNOR2_X1 U382 ( .A(n526), .B(KEYINPUT68), .ZN(n379) );
  XNOR2_X2 U383 ( .A(n537), .B(KEYINPUT102), .ZN(n577) );
  XNOR2_X2 U384 ( .A(n394), .B(n340), .ZN(n548) );
  NOR2_X4 U385 ( .A1(n684), .A2(n615), .ZN(n689) );
  XNOR2_X1 U386 ( .A(n596), .B(KEYINPUT79), .ZN(n361) );
  NAND2_X1 U387 ( .A1(n356), .A2(n355), .ZN(n354) );
  NAND2_X1 U388 ( .A1(n430), .A2(G902), .ZN(n355) );
  NAND2_X1 U389 ( .A1(n702), .A2(n430), .ZN(n356) );
  XOR2_X1 U390 ( .A(KEYINPUT4), .B(G137), .Z(n526) );
  XNOR2_X1 U391 ( .A(G146), .B(G125), .ZN(n460) );
  XNOR2_X1 U392 ( .A(n360), .B(n598), .ZN(n412) );
  XNOR2_X1 U393 ( .A(n444), .B(n445), .ZN(n346) );
  NAND2_X1 U394 ( .A1(n726), .A2(G227), .ZN(n445) );
  XNOR2_X1 U395 ( .A(n529), .B(n531), .ZN(n444) );
  XNOR2_X1 U396 ( .A(n446), .B(KEYINPUT67), .ZN(n530) );
  INV_X1 U397 ( .A(G140), .ZN(n446) );
  XNOR2_X1 U398 ( .A(KEYINPUT4), .B(KEYINPUT75), .ZN(n482) );
  XOR2_X1 U399 ( .A(KEYINPUT87), .B(KEYINPUT18), .Z(n483) );
  XNOR2_X1 U400 ( .A(n485), .B(n409), .ZN(n408) );
  INV_X1 U401 ( .A(KEYINPUT17), .ZN(n409) );
  INV_X1 U402 ( .A(n460), .ZN(n486) );
  XNOR2_X1 U403 ( .A(n414), .B(G128), .ZN(n509) );
  INV_X1 U404 ( .A(G143), .ZN(n414) );
  INV_X1 U405 ( .A(KEYINPUT44), .ZN(n384) );
  INV_X1 U406 ( .A(KEYINPUT19), .ZN(n493) );
  AND2_X1 U407 ( .A1(n348), .A2(n347), .ZN(n661) );
  AND2_X1 U408 ( .A1(n350), .A2(n565), .ZN(n348) );
  INV_X1 U409 ( .A(n354), .ZN(n347) );
  INV_X1 U410 ( .A(G146), .ZN(n531) );
  XOR2_X1 U411 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n522) );
  XNOR2_X1 U412 ( .A(n532), .B(n432), .ZN(n431) );
  XNOR2_X1 U413 ( .A(n433), .B(KEYINPUT16), .ZN(n432) );
  INV_X1 U414 ( .A(G122), .ZN(n433) );
  XNOR2_X1 U415 ( .A(n509), .B(n413), .ZN(n527) );
  INV_X1 U416 ( .A(G134), .ZN(n413) );
  NOR2_X1 U417 ( .A1(n646), .A2(n612), .ZN(n613) );
  AND2_X1 U418 ( .A1(n438), .A2(n336), .ZN(n437) );
  XNOR2_X1 U419 ( .A(G469), .B(KEYINPUT70), .ZN(n447) );
  OR2_X1 U420 ( .A1(n694), .A2(G902), .ZN(n448) );
  NOR2_X1 U421 ( .A1(n371), .A2(G902), .ZN(n416) );
  OR2_X1 U422 ( .A1(n354), .A2(n349), .ZN(n664) );
  INV_X1 U423 ( .A(n350), .ZN(n349) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n469) );
  INV_X1 U425 ( .A(G101), .ZN(n529) );
  XNOR2_X1 U426 ( .A(n654), .B(KEYINPUT80), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n380), .B(G131), .ZN(n525) );
  INV_X1 U428 ( .A(KEYINPUT66), .ZN(n380) );
  XOR2_X1 U429 ( .A(G140), .B(KEYINPUT11), .Z(n458) );
  NAND2_X1 U430 ( .A1(n462), .A2(n461), .ZN(n429) );
  XNOR2_X1 U431 ( .A(n525), .B(KEYINPUT12), .ZN(n368) );
  XNOR2_X1 U432 ( .A(G113), .B(G143), .ZN(n455) );
  XOR2_X1 U433 ( .A(G104), .B(G122), .Z(n456) );
  XNOR2_X1 U434 ( .A(n584), .B(KEYINPUT46), .ZN(n427) );
  NOR2_X1 U435 ( .A1(n730), .A2(n733), .ZN(n584) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n495) );
  NAND2_X1 U437 ( .A1(n439), .A2(KEYINPUT34), .ZN(n438) );
  INV_X1 U438 ( .A(n558), .ZN(n439) );
  INV_X1 U439 ( .A(KEYINPUT0), .ZN(n393) );
  OR2_X1 U440 ( .A1(n351), .A2(n702), .ZN(n350) );
  NAND2_X1 U441 ( .A1(n353), .A2(n352), .ZN(n351) );
  INV_X1 U442 ( .A(G902), .ZN(n352) );
  INV_X1 U443 ( .A(n430), .ZN(n353) );
  XNOR2_X1 U444 ( .A(n359), .B(KEYINPUT24), .ZN(n358) );
  XNOR2_X1 U445 ( .A(KEYINPUT82), .B(KEYINPUT23), .ZN(n359) );
  XNOR2_X1 U446 ( .A(G119), .B(G137), .ZN(n357) );
  XNOR2_X1 U447 ( .A(n429), .B(n428), .ZN(n716) );
  INV_X1 U448 ( .A(n530), .ZN(n428) );
  XNOR2_X1 U449 ( .A(G128), .B(G110), .ZN(n464) );
  XOR2_X1 U450 ( .A(KEYINPUT93), .B(KEYINPUT71), .Z(n465) );
  XNOR2_X1 U451 ( .A(G116), .B(G122), .ZN(n513) );
  XNOR2_X1 U452 ( .A(n369), .B(n367), .ZN(n506) );
  XNOR2_X1 U453 ( .A(n463), .B(n370), .ZN(n369) );
  XNOR2_X1 U454 ( .A(n429), .B(n368), .ZN(n367) );
  XNOR2_X1 U455 ( .A(n457), .B(n458), .ZN(n370) );
  XNOR2_X1 U456 ( .A(n535), .B(n715), .ZN(n694) );
  XNOR2_X1 U457 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U458 ( .A(n346), .B(n530), .ZN(n534) );
  XNOR2_X1 U459 ( .A(n484), .B(n408), .ZN(n487) );
  INV_X1 U460 ( .A(KEYINPUT45), .ZN(n434) );
  XNOR2_X1 U461 ( .A(n382), .B(KEYINPUT101), .ZN(n381) );
  AND2_X1 U462 ( .A1(n648), .A2(n582), .ZN(n583) );
  NAND2_X1 U463 ( .A1(n636), .A2(n417), .ZN(n607) );
  AND2_X1 U464 ( .A1(n600), .A2(n418), .ZN(n417) );
  NOR2_X1 U465 ( .A1(n601), .A2(n419), .ZN(n418) );
  NAND2_X1 U466 ( .A1(n602), .A2(n649), .ZN(n419) );
  AND2_X1 U467 ( .A1(n661), .A2(n581), .ZN(n589) );
  XNOR2_X1 U468 ( .A(n335), .B(n715), .ZN(n371) );
  XNOR2_X1 U469 ( .A(n422), .B(n420), .ZN(n699) );
  XNOR2_X1 U470 ( .A(n512), .B(n421), .ZN(n420) );
  XNOR2_X1 U471 ( .A(n515), .B(n527), .ZN(n422) );
  XNOR2_X1 U472 ( .A(n513), .B(KEYINPUT7), .ZN(n421) );
  NAND2_X1 U473 ( .A1(n375), .A2(n372), .ZN(n730) );
  NAND2_X1 U474 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X1 U475 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U476 ( .A1(n599), .A2(n378), .ZN(n373) );
  XNOR2_X1 U477 ( .A(n547), .B(n546), .ZN(n731) );
  INV_X1 U478 ( .A(n586), .ZN(n365) );
  OR2_X1 U479 ( .A1(n577), .A2(n397), .ZN(n396) );
  INV_X1 U480 ( .A(n664), .ZN(n397) );
  NOR2_X1 U481 ( .A1(n664), .A2(n550), .ZN(n619) );
  XNOR2_X1 U482 ( .A(n549), .B(KEYINPUT83), .ZN(n550) );
  NOR2_X1 U483 ( .A1(n548), .A2(n406), .ZN(n549) );
  OR2_X1 U484 ( .A1(n600), .A2(n407), .ZN(n406) );
  XNOR2_X1 U485 ( .A(n701), .B(n702), .ZN(n395) );
  INV_X1 U486 ( .A(KEYINPUT120), .ZN(n401) );
  INV_X1 U487 ( .A(KEYINPUT56), .ZN(n398) );
  XNOR2_X1 U488 ( .A(n494), .B(n493), .ZN(n585) );
  XOR2_X1 U489 ( .A(n492), .B(n491), .Z(n334) );
  XOR2_X1 U490 ( .A(n519), .B(n524), .Z(n335) );
  XOR2_X1 U491 ( .A(n588), .B(KEYINPUT76), .Z(n336) );
  XOR2_X1 U492 ( .A(n587), .B(KEYINPUT73), .Z(n337) );
  INV_X1 U493 ( .A(n606), .ZN(n407) );
  NOR2_X1 U494 ( .A1(n503), .A2(n393), .ZN(n338) );
  NAND2_X1 U495 ( .A1(n664), .A2(n407), .ZN(n339) );
  INV_X1 U496 ( .A(KEYINPUT34), .ZN(n443) );
  XOR2_X1 U497 ( .A(n518), .B(KEYINPUT64), .Z(n340) );
  XNOR2_X1 U498 ( .A(n696), .B(n695), .ZN(n341) );
  XNOR2_X1 U499 ( .A(n506), .B(KEYINPUT59), .ZN(n342) );
  XOR2_X1 U500 ( .A(n371), .B(n618), .Z(n343) );
  XOR2_X1 U501 ( .A(n692), .B(n691), .Z(n344) );
  NOR2_X1 U502 ( .A1(G952), .A2(n726), .ZN(n703) );
  INV_X1 U503 ( .A(n703), .ZN(n452) );
  XOR2_X1 U504 ( .A(n617), .B(KEYINPUT65), .Z(n345) );
  NAND2_X1 U505 ( .A1(n558), .A2(n517), .ZN(n394) );
  NAND2_X1 U506 ( .A1(n440), .A2(n437), .ZN(n436) );
  NAND2_X1 U507 ( .A1(n337), .A2(n364), .ZN(n363) );
  INV_X1 U508 ( .A(n633), .ZN(n364) );
  NOR2_X1 U509 ( .A1(n366), .A2(KEYINPUT47), .ZN(n587) );
  NOR2_X1 U510 ( .A1(n563), .A2(n366), .ZN(n564) );
  INV_X1 U511 ( .A(n611), .ZN(n374) );
  NAND2_X1 U512 ( .A1(n599), .A2(n378), .ZN(n376) );
  NAND2_X1 U513 ( .A1(n611), .A2(n378), .ZN(n377) );
  INV_X1 U514 ( .A(KEYINPUT40), .ZN(n378) );
  NAND2_X1 U515 ( .A1(n383), .A2(n381), .ZN(n435) );
  OR2_X1 U516 ( .A1(n564), .A2(n619), .ZN(n382) );
  XNOR2_X1 U517 ( .A(n385), .B(n384), .ZN(n383) );
  NAND2_X1 U518 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U519 ( .A(n731), .ZN(n386) );
  XNOR2_X1 U520 ( .A(n541), .B(KEYINPUT84), .ZN(n387) );
  NAND2_X1 U521 ( .A1(n585), .A2(n393), .ZN(n392) );
  INV_X1 U522 ( .A(n585), .ZN(n389) );
  NOR2_X2 U523 ( .A1(n707), .A2(n724), .ZN(n614) );
  XNOR2_X2 U524 ( .A(n614), .B(KEYINPUT2), .ZN(n684) );
  XNOR2_X1 U525 ( .A(n540), .B(KEYINPUT32), .ZN(n732) );
  NOR2_X1 U526 ( .A1(n395), .A2(n703), .ZN(G66) );
  OR2_X2 U527 ( .A1(n548), .A2(n396), .ZN(n536) );
  XNOR2_X1 U528 ( .A(n399), .B(n398), .ZN(G51) );
  NAND2_X1 U529 ( .A1(n403), .A2(n452), .ZN(n399) );
  XNOR2_X1 U530 ( .A(n400), .B(n345), .ZN(G60) );
  NAND2_X1 U531 ( .A1(n405), .A2(n452), .ZN(n400) );
  XNOR2_X1 U532 ( .A(n402), .B(n401), .ZN(G54) );
  NAND2_X1 U533 ( .A1(n404), .A2(n452), .ZN(n402) );
  XNOR2_X1 U534 ( .A(n693), .B(n344), .ZN(n403) );
  XNOR2_X1 U535 ( .A(n697), .B(n341), .ZN(n404) );
  NAND2_X1 U536 ( .A1(n412), .A2(n411), .ZN(n410) );
  XNOR2_X1 U537 ( .A(n410), .B(KEYINPUT69), .ZN(n426) );
  XNOR2_X2 U538 ( .A(n415), .B(n527), .ZN(n715) );
  XNOR2_X1 U539 ( .A(n616), .B(n342), .ZN(n405) );
  NAND2_X1 U540 ( .A1(n690), .A2(n615), .ZN(n450) );
  XNOR2_X1 U541 ( .A(n489), .B(n488), .ZN(n690) );
  INV_X1 U542 ( .A(n642), .ZN(n411) );
  XNOR2_X2 U543 ( .A(n416), .B(n528), .ZN(n537) );
  NAND2_X1 U544 ( .A1(n423), .A2(n613), .ZN(n724) );
  XNOR2_X1 U545 ( .A(n425), .B(n424), .ZN(n423) );
  INV_X1 U546 ( .A(KEYINPUT48), .ZN(n424) );
  NAND2_X1 U547 ( .A1(n427), .A2(n426), .ZN(n425) );
  NAND2_X1 U548 ( .A1(n659), .A2(n441), .ZN(n440) );
  AND2_X1 U549 ( .A1(n558), .A2(n443), .ZN(n441) );
  NOR2_X1 U550 ( .A1(n659), .A2(n443), .ZN(n442) );
  XNOR2_X2 U551 ( .A(n545), .B(KEYINPUT33), .ZN(n659) );
  XNOR2_X2 U552 ( .A(n448), .B(n447), .ZN(n581) );
  XNOR2_X2 U553 ( .A(n449), .B(n480), .ZN(n519) );
  NAND2_X1 U554 ( .A1(n610), .A2(n649), .ZN(n494) );
  XNOR2_X2 U555 ( .A(n450), .B(n334), .ZN(n610) );
  NAND2_X1 U556 ( .A1(n529), .A2(KEYINPUT3), .ZN(n477) );
  XNOR2_X1 U557 ( .A(n451), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U558 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n454), .B(n343), .ZN(n453) );
  NAND2_X1 U560 ( .A1(n689), .A2(G472), .ZN(n454) );
  NOR2_X2 U561 ( .A1(n536), .A2(n407), .ZN(n627) );
  INV_X1 U562 ( .A(KEYINPUT72), .ZN(n598) );
  XNOR2_X1 U563 ( .A(n523), .B(n531), .ZN(n524) );
  INV_X1 U564 ( .A(G472), .ZN(n528) );
  INV_X1 U565 ( .A(n645), .ZN(n612) );
  XOR2_X1 U566 ( .A(n538), .B(KEYINPUT100), .Z(n600) );
  XNOR2_X1 U567 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U568 ( .A(n456), .B(n455), .ZN(n463) );
  NAND2_X1 U569 ( .A1(G214), .A2(n520), .ZN(n457) );
  INV_X1 U570 ( .A(KEYINPUT10), .ZN(n459) );
  NAND2_X1 U571 ( .A1(n486), .A2(n459), .ZN(n462) );
  NAND2_X1 U572 ( .A1(n460), .A2(KEYINPUT10), .ZN(n461) );
  XNOR2_X1 U573 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n716), .B(n466), .ZN(n471) );
  NAND2_X1 U575 ( .A1(G234), .A2(n726), .ZN(n467) );
  XOR2_X1 U576 ( .A(KEYINPUT8), .B(n467), .Z(n514) );
  NAND2_X1 U577 ( .A1(n514), .A2(G221), .ZN(n468) );
  XNOR2_X1 U578 ( .A(G902), .B(KEYINPUT15), .ZN(n615) );
  NAND2_X1 U579 ( .A1(n615), .A2(G234), .ZN(n473) );
  XNOR2_X1 U580 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n473), .B(n472), .ZN(n504) );
  NAND2_X1 U582 ( .A1(G217), .A2(n504), .ZN(n474) );
  OR2_X1 U583 ( .A1(G237), .A2(G902), .ZN(n490) );
  NAND2_X1 U584 ( .A1(G214), .A2(n490), .ZN(n649) );
  INV_X1 U585 ( .A(KEYINPUT3), .ZN(n476) );
  NAND2_X1 U586 ( .A1(n476), .A2(G101), .ZN(n478) );
  NAND2_X1 U587 ( .A1(n478), .A2(n477), .ZN(n480) );
  XNOR2_X2 U588 ( .A(G119), .B(KEYINPUT86), .ZN(n481) );
  XNOR2_X1 U589 ( .A(n710), .B(n509), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U591 ( .A1(G224), .A2(n726), .ZN(n485) );
  XOR2_X1 U592 ( .A(n487), .B(n486), .Z(n488) );
  XOR2_X1 U593 ( .A(KEYINPUT77), .B(KEYINPUT88), .Z(n492) );
  NAND2_X1 U594 ( .A1(G210), .A2(n490), .ZN(n491) );
  XNOR2_X1 U595 ( .A(n495), .B(KEYINPUT14), .ZN(n497) );
  NAND2_X1 U596 ( .A1(n497), .A2(G952), .ZN(n496) );
  XOR2_X1 U597 ( .A(KEYINPUT89), .B(n496), .Z(n679) );
  NOR2_X1 U598 ( .A1(G953), .A2(n679), .ZN(n569) );
  NAND2_X1 U599 ( .A1(G902), .A2(n497), .ZN(n498) );
  XOR2_X1 U600 ( .A(KEYINPUT90), .B(n498), .Z(n499) );
  NAND2_X1 U601 ( .A1(G953), .A2(n499), .ZN(n566) );
  NOR2_X1 U602 ( .A1(G898), .A2(n566), .ZN(n500) );
  XOR2_X1 U603 ( .A(KEYINPUT91), .B(n500), .Z(n501) );
  NOR2_X1 U604 ( .A1(n569), .A2(n501), .ZN(n502) );
  XNOR2_X1 U605 ( .A(n502), .B(KEYINPUT92), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n504), .A2(G221), .ZN(n505) );
  XOR2_X1 U607 ( .A(KEYINPUT21), .B(n505), .Z(n565) );
  XNOR2_X1 U608 ( .A(KEYINPUT13), .B(G475), .ZN(n508) );
  NOR2_X1 U609 ( .A1(G902), .A2(n506), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n508), .B(n507), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n511) );
  XNOR2_X1 U612 ( .A(G107), .B(KEYINPUT9), .ZN(n510) );
  XNOR2_X1 U613 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U614 ( .A1(G217), .A2(n514), .ZN(n515) );
  NOR2_X1 U615 ( .A1(G902), .A2(n699), .ZN(n516) );
  XOR2_X1 U616 ( .A(G478), .B(n516), .Z(n553) );
  NOR2_X1 U617 ( .A1(n551), .A2(n553), .ZN(n574) );
  AND2_X1 U618 ( .A1(n565), .A2(n574), .ZN(n517) );
  INV_X1 U619 ( .A(KEYINPUT22), .ZN(n518) );
  NAND2_X1 U620 ( .A1(n520), .A2(G210), .ZN(n521) );
  XNOR2_X1 U621 ( .A(n522), .B(n521), .ZN(n523) );
  INV_X1 U622 ( .A(n532), .ZN(n533) );
  XNOR2_X1 U623 ( .A(KEYINPUT1), .B(n581), .ZN(n542) );
  INV_X1 U624 ( .A(n542), .ZN(n606) );
  XNOR2_X1 U625 ( .A(n537), .B(KEYINPUT6), .ZN(n538) );
  OR2_X1 U626 ( .A1(n600), .A2(n339), .ZN(n539) );
  NAND2_X1 U627 ( .A1(n551), .A2(n553), .ZN(n588) );
  INV_X1 U628 ( .A(n565), .ZN(n663) );
  NAND2_X1 U629 ( .A1(n661), .A2(n542), .ZN(n543) );
  XNOR2_X2 U630 ( .A(n543), .B(KEYINPUT74), .ZN(n555) );
  XNOR2_X1 U631 ( .A(n555), .B(KEYINPUT103), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n544), .A2(n600), .ZN(n545) );
  INV_X1 U633 ( .A(KEYINPUT35), .ZN(n546) );
  INV_X1 U634 ( .A(n551), .ZN(n552) );
  OR2_X1 U635 ( .A1(n552), .A2(n553), .ZN(n599) );
  NAND2_X1 U636 ( .A1(n553), .A2(n552), .ZN(n628) );
  AND2_X1 U637 ( .A1(n599), .A2(n628), .ZN(n654) );
  XOR2_X1 U638 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n557) );
  INV_X1 U639 ( .A(n537), .ZN(n554) );
  NOR2_X1 U640 ( .A1(n555), .A2(n554), .ZN(n671) );
  NAND2_X1 U641 ( .A1(n671), .A2(n558), .ZN(n556) );
  XNOR2_X1 U642 ( .A(n557), .B(n556), .ZN(n640) );
  INV_X1 U643 ( .A(n581), .ZN(n560) );
  NAND2_X1 U644 ( .A1(n661), .A2(n558), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U646 ( .A(n561), .B(KEYINPUT95), .ZN(n562) );
  NOR2_X1 U647 ( .A1(n537), .A2(n562), .ZN(n622) );
  NOR2_X1 U648 ( .A1(n640), .A2(n622), .ZN(n563) );
  NAND2_X1 U649 ( .A1(n664), .A2(n565), .ZN(n601) );
  NOR2_X1 U650 ( .A1(G900), .A2(n566), .ZN(n567) );
  XOR2_X1 U651 ( .A(KEYINPUT105), .B(n567), .Z(n568) );
  NOR2_X1 U652 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U653 ( .A(KEYINPUT78), .B(n570), .Z(n602) );
  NAND2_X1 U654 ( .A1(n602), .A2(n577), .ZN(n571) );
  XNOR2_X1 U655 ( .A(n572), .B(KEYINPUT28), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n573), .A2(n581), .ZN(n586) );
  INV_X1 U657 ( .A(n610), .ZN(n603) );
  XNOR2_X1 U658 ( .A(n603), .B(KEYINPUT38), .ZN(n648) );
  NAND2_X1 U659 ( .A1(n649), .A2(n648), .ZN(n653) );
  INV_X1 U660 ( .A(n574), .ZN(n651) );
  NOR2_X1 U661 ( .A1(n653), .A2(n651), .ZN(n575) );
  XNOR2_X1 U662 ( .A(KEYINPUT41), .B(n575), .ZN(n680) );
  NOR2_X1 U663 ( .A1(n586), .A2(n680), .ZN(n576) );
  XNOR2_X1 U664 ( .A(n576), .B(KEYINPUT42), .ZN(n733) );
  NAND2_X1 U665 ( .A1(n577), .A2(n649), .ZN(n579) );
  XOR2_X1 U666 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n578) );
  XNOR2_X1 U667 ( .A(n579), .B(n578), .ZN(n580) );
  AND2_X1 U668 ( .A1(n580), .A2(n602), .ZN(n593) );
  AND2_X1 U669 ( .A1(n593), .A2(n589), .ZN(n582) );
  INV_X1 U670 ( .A(n588), .ZN(n591) );
  AND2_X1 U671 ( .A1(n610), .A2(n589), .ZN(n590) );
  AND2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U673 ( .A(n632), .B(KEYINPUT81), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n654), .A2(KEYINPUT47), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U676 ( .A1(KEYINPUT47), .A2(n633), .ZN(n597) );
  XNOR2_X1 U677 ( .A(KEYINPUT104), .B(n599), .ZN(n634) );
  INV_X1 U678 ( .A(n634), .ZN(n636) );
  XOR2_X1 U679 ( .A(KEYINPUT36), .B(n604), .Z(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n642) );
  NOR2_X1 U681 ( .A1(n407), .A2(n607), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT43), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n646) );
  OR2_X1 U684 ( .A1(n628), .A2(n611), .ZN(n645) );
  NAND2_X1 U685 ( .A1(n689), .A2(G475), .ZN(n616) );
  INV_X1 U686 ( .A(KEYINPUT60), .ZN(n617) );
  XOR2_X1 U687 ( .A(KEYINPUT62), .B(KEYINPUT85), .Z(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(G101), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(KEYINPUT107), .ZN(G3) );
  NAND2_X1 U690 ( .A1(n636), .A2(n622), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n621), .B(G104), .ZN(G6) );
  XNOR2_X1 U692 ( .A(G107), .B(KEYINPUT27), .ZN(n626) );
  XOR2_X1 U693 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n624) );
  INV_X1 U694 ( .A(n628), .ZN(n639) );
  NAND2_X1 U695 ( .A1(n622), .A2(n639), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(G9) );
  XOR2_X1 U698 ( .A(n627), .B(G110), .Z(G12) );
  NOR2_X1 U699 ( .A1(n628), .A2(n633), .ZN(n630) );
  XNOR2_X1 U700 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(n631) );
  XOR2_X1 U702 ( .A(G128), .B(n631), .Z(G30) );
  XOR2_X1 U703 ( .A(n632), .B(G143), .Z(G45) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(G146), .B(n635), .Z(G48) );
  NAND2_X1 U706 ( .A1(n636), .A2(n640), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT110), .ZN(n638) );
  XNOR2_X1 U708 ( .A(G113), .B(n638), .ZN(G15) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(G116), .ZN(G18) );
  XOR2_X1 U711 ( .A(KEYINPUT111), .B(KEYINPUT37), .Z(n644) );
  XNOR2_X1 U712 ( .A(n642), .B(G125), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n645), .ZN(G36) );
  XOR2_X1 U715 ( .A(G140), .B(n646), .Z(n647) );
  XNOR2_X1 U716 ( .A(KEYINPUT112), .B(n647), .ZN(G42) );
  NOR2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U719 ( .A(KEYINPUT115), .B(n652), .Z(n657) );
  NOR2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U721 ( .A(KEYINPUT116), .B(n655), .ZN(n656) );
  NOR2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U723 ( .A(KEYINPUT117), .B(n658), .ZN(n660) );
  NAND2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n676) );
  NOR2_X1 U725 ( .A1(n407), .A2(n661), .ZN(n662) );
  XOR2_X1 U726 ( .A(KEYINPUT50), .B(n662), .Z(n668) );
  NAND2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U728 ( .A(n665), .B(KEYINPUT49), .ZN(n666) );
  XNOR2_X1 U729 ( .A(KEYINPUT113), .B(n666), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U731 ( .A1(n537), .A2(n669), .ZN(n670) );
  NOR2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U733 ( .A(KEYINPUT51), .B(n672), .Z(n673) );
  NOR2_X1 U734 ( .A1(n680), .A2(n673), .ZN(n674) );
  XOR2_X1 U735 ( .A(KEYINPUT114), .B(n674), .Z(n675) );
  NAND2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U737 ( .A(KEYINPUT52), .B(n677), .Z(n678) );
  NOR2_X1 U738 ( .A1(n679), .A2(n678), .ZN(n683) );
  INV_X1 U739 ( .A(n659), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U743 ( .A(KEYINPUT118), .B(n686), .ZN(n687) );
  NOR2_X1 U744 ( .A1(n687), .A2(G953), .ZN(n688) );
  XNOR2_X1 U745 ( .A(n688), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U746 ( .A1(n689), .A2(G210), .ZN(n693) );
  INV_X1 U747 ( .A(n690), .ZN(n692) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n691) );
  NAND2_X1 U749 ( .A1(n689), .A2(G469), .ZN(n697) );
  XOR2_X1 U750 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  XNOR2_X1 U751 ( .A(n694), .B(KEYINPUT119), .ZN(n695) );
  NAND2_X1 U752 ( .A1(G478), .A2(n689), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n703), .A2(n700), .ZN(G63) );
  NAND2_X1 U755 ( .A1(G217), .A2(n689), .ZN(n701) );
  INV_X1 U756 ( .A(G898), .ZN(n706) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n704) );
  XOR2_X1 U758 ( .A(KEYINPUT61), .B(n704), .Z(n705) );
  NOR2_X1 U759 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U760 ( .A1(G953), .A2(n707), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U762 ( .A1(G898), .A2(n726), .ZN(n712) );
  XOR2_X1 U763 ( .A(n710), .B(KEYINPUT121), .Z(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U765 ( .A(n714), .B(n713), .Z(G69) );
  XNOR2_X1 U766 ( .A(G227), .B(KEYINPUT123), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(n722) );
  INV_X1 U768 ( .A(n722), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(n719) );
  NAND2_X1 U770 ( .A1(G900), .A2(n719), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n720), .B(KEYINPUT124), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n721), .A2(G953), .ZN(n728) );
  XNOR2_X1 U773 ( .A(n722), .B(KEYINPUT122), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(G72) );
  XOR2_X1 U777 ( .A(G131), .B(KEYINPUT126), .Z(n729) );
  XNOR2_X1 U778 ( .A(n730), .B(n729), .ZN(G33) );
  XOR2_X1 U779 ( .A(G122), .B(n731), .Z(G24) );
  XOR2_X1 U780 ( .A(n732), .B(G119), .Z(G21) );
  XNOR2_X1 U781 ( .A(G137), .B(KEYINPUT125), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(n733), .ZN(G39) );
endmodule

