//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT11), .B(G169gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G43gat), .A2(G50gat), .ZN(new_n215));
  AND2_X1   g014(.A1(G43gat), .A2(G50gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(KEYINPUT15), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n220));
  AND4_X1   g019(.A1(new_n212), .A2(new_n210), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT15), .B1(new_n216), .B2(new_n215), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(G43gat), .A2(G50gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT89), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n225), .A2(new_n230), .A3(new_n226), .A4(new_n227), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n221), .A2(new_n222), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G22gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G15gat), .ZN(new_n234));
  INV_X1    g033(.A(G15gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G22gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G1gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(KEYINPUT16), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n234), .A3(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G8gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(KEYINPUT91), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n240), .A2(new_n234), .A3(new_n236), .A4(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT92), .B(G8gat), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n244), .A2(new_n239), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n217), .A2(new_n232), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n248), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n229), .A2(new_n231), .ZN(new_n256));
  AND3_X1   g055(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(new_n222), .A3(new_n212), .A4(new_n210), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n255), .B(new_n217), .C1(new_n256), .C2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n255), .B1(new_n232), .B2(new_n217), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n217), .B1(new_n256), .B2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT17), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n261), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT93), .A3(new_n254), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n252), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(new_n251), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT97), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n232), .A2(new_n243), .A3(new_n248), .A4(new_n217), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n249), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(new_n274), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n271), .A2(KEYINPUT18), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT95), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n207), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT18), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n271), .B2(KEYINPUT94), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n249), .B1(G229gat), .B2(G233gat), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT93), .B1(new_n269), .B2(new_n254), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n265), .B(new_n253), .C1(new_n268), .C2(new_n261), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT94), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n279), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT18), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n278), .A2(new_n273), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT18), .B1(new_n287), .B2(new_n288), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n271), .A2(KEYINPUT94), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n206), .B1(new_n294), .B2(KEYINPUT95), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G197gat), .B(G204gat), .ZN(new_n302));
  INV_X1    g101(.A(G211gat), .ZN(new_n303));
  INV_X1    g102(.A(G218gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(KEYINPUT22), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT74), .ZN(new_n309));
  INV_X1    g108(.A(G226gat), .ZN(new_n310));
  INV_X1    g109(.A(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n314), .A2(KEYINPUT25), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT64), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT64), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT65), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n318), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n314), .A2(new_n317), .A3(new_n316), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n325), .B1(new_n319), .B2(new_n320), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n327), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT25), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n313), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  INV_X1    g133(.A(G169gat), .ZN(new_n335));
  INV_X1    g134(.A(G176gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT27), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G183gat), .ZN(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT28), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT27), .B(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n346), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n334), .B2(new_n339), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n329), .A2(new_n333), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n312), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n312), .ZN(new_n357));
  INV_X1    g156(.A(new_n319), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT64), .B(KEYINPUT24), .ZN(new_n359));
  INV_X1    g158(.A(new_n325), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n327), .B(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT25), .B(new_n330), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n331), .A2(new_n327), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n314), .A2(new_n317), .A3(new_n316), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n353), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n370), .A2(new_n341), .A3(new_n351), .A4(new_n348), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n357), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n309), .B1(new_n356), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT75), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n312), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n369), .B2(new_n371), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n308), .B(new_n379), .C1(new_n380), .C2(new_n312), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(new_n381), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n377), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT30), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT76), .B1(new_n383), .B2(new_n377), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n388));
  AOI211_X1 g187(.A(new_n388), .B(new_n378), .C1(new_n373), .C2(new_n381), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n390), .B2(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(G113gat), .ZN(new_n392));
  INV_X1    g191(.A(G120gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT1), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G113gat), .A2(G120gat), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G127gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n398));
  INV_X1    g197(.A(G134gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G127gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT68), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n404), .A2(KEYINPUT67), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(KEYINPUT67), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n400), .B(new_n398), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n396), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT69), .B(G113gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(new_n393), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n397), .A2(G134gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n400), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n416));
  INV_X1    g215(.A(G148gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(G141gat), .ZN(new_n418));
  INV_X1    g217(.A(G141gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(G148gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT77), .B1(new_n417), .B2(G141gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n419), .A3(G148gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n417), .A2(G141gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n422), .B2(KEYINPUT2), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT3), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n421), .A2(new_n424), .B1(new_n430), .B2(new_n431), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n439), .A3(KEYINPUT3), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n415), .A2(new_n435), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n407), .A2(new_n403), .ZN(new_n443));
  INV_X1    g242(.A(new_n396), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n413), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n436), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n447), .A2(KEYINPUT4), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(KEYINPUT4), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n441), .B(new_n442), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451));
  INV_X1    g250(.A(new_n442), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n408), .A2(new_n433), .A3(new_n413), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n436), .B1(new_n445), .B2(new_n446), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n455), .B2(KEYINPUT5), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n433), .B1(new_n408), .B2(new_n413), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n442), .B1(new_n447), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT5), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n458), .A2(KEYINPUT80), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n450), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  XOR2_X1   g261(.A(G1gat), .B(G29gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G57gat), .B(G85gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n447), .B(KEYINPUT4), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(new_n459), .A3(new_n442), .A4(new_n441), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n461), .A2(new_n462), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n461), .A2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n461), .B2(new_n470), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n468), .A3(new_n470), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(KEYINPUT82), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n391), .B(new_n476), .C1(new_n479), .C2(KEYINPUT6), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n478), .A2(KEYINPUT82), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT6), .B1(new_n482), .B2(new_n475), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n391), .A4(new_n476), .ZN(new_n486));
  INV_X1    g285(.A(new_n307), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n306), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n355), .A3(new_n433), .ZN(new_n489));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(new_n434), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n438), .A2(new_n355), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n488), .B(KEYINPUT74), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n496));
  INV_X1    g295(.A(new_n437), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n433), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n308), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT85), .B(G22gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G78gat), .B(G106gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(new_n224), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT86), .B1(new_n501), .B2(new_n233), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(G22gat), .C1(new_n495), .C2(new_n500), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n501), .B2(new_n502), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n503), .A2(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n481), .A2(new_n486), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n354), .B(new_n414), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n515), .A2(KEYINPUT72), .B1(G227gat), .B2(G233gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(KEYINPUT72), .B2(new_n515), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT34), .ZN(new_n520));
  NAND2_X1  g319(.A1(G227gat), .A2(G233gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT32), .B1(new_n515), .B2(new_n521), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n515), .B2(new_n521), .ZN(new_n527));
  XOR2_X1   g326(.A(G15gat), .B(G43gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT70), .ZN(new_n529));
  XOR2_X1   g328(.A(G71gat), .B(G99gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  OAI221_X1 g332(.A(KEYINPUT32), .B1(new_n526), .B2(new_n531), .C1(new_n515), .C2(new_n521), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n519), .A2(new_n523), .A3(new_n534), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n514), .A2(KEYINPUT87), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT87), .B1(new_n514), .B2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n384), .A2(new_n388), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n378), .B1(new_n373), .B2(new_n381), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n385), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n386), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n447), .A2(new_n457), .A3(new_n442), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT39), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n469), .A2(new_n441), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(new_n452), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT39), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n556), .A3(new_n452), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT40), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n467), .B1(KEYINPUT88), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n555), .A2(new_n557), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n559), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n562), .A2(new_n554), .B1(KEYINPUT88), .B2(new_n558), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n550), .A2(new_n475), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n503), .A2(new_n507), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n511), .A2(new_n512), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n477), .B1(new_n472), .B2(new_n471), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n483), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n377), .B1(new_n383), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n570), .B2(new_n383), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT38), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n356), .A2(new_n372), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n494), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n575), .B(KEYINPUT37), .C1(new_n308), .C2(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n390), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n564), .B(new_n567), .C1(new_n569), .C2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n543), .A2(new_n544), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n536), .A3(new_n537), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n583), .A2(new_n480), .A3(KEYINPUT35), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n538), .A2(new_n513), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n485), .B1(new_n569), .B2(new_n391), .ZN(new_n586));
  NOR4_X1   g385(.A1(new_n483), .A2(new_n550), .A3(new_n568), .A4(KEYINPUT83), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n584), .B1(new_n588), .B2(KEYINPUT35), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n301), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT7), .ZN(new_n593));
  OR2_X1    g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT101), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n603), .A2(new_n593), .A3(new_n596), .A4(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n267), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT41), .ZN(new_n609));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n268), .B2(new_n261), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT102), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n609), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT100), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  OAI21_X1  g420(.A(new_n615), .B1(new_n611), .B2(new_n612), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(KEYINPUT103), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n617), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n613), .A2(KEYINPUT103), .A3(new_n616), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G57gat), .B(G64gat), .Z(new_n632));
  NAND2_X1  g431(.A1(G71gat), .A2(G78gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT9), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n633), .A2(new_n638), .B1(new_n635), .B2(KEYINPUT98), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n633), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n637), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n632), .B(new_n635), .C1(new_n642), .C2(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT21), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(G127gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n253), .B1(KEYINPUT21), .B2(new_n644), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT99), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(G127gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n651), .B1(new_n655), .B2(new_n648), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G155gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G183gat), .B(G211gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n654), .B2(new_n656), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n596), .A2(new_n599), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n603), .B1(new_n665), .B2(new_n593), .ZN(new_n666));
  AND4_X1   g465(.A1(new_n603), .A2(new_n593), .A3(new_n596), .A4(new_n599), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n644), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n605), .A2(new_n640), .A3(new_n606), .A4(new_n643), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n644), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G230gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n311), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n668), .B2(new_n670), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G120gat), .B(G148gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  NAND3_X1  g481(.A1(new_n677), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n675), .B1(new_n671), .B2(new_n672), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n678), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n631), .A2(new_n664), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n591), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n569), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n238), .ZN(G1324gat));
  XOR2_X1   g494(.A(KEYINPUT16), .B(G8gat), .Z(new_n696));
  NAND4_X1  g495(.A1(new_n591), .A2(new_n550), .A3(new_n688), .A4(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G8gat), .B1(new_n689), .B2(new_n391), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n697), .ZN(new_n699));
  MUX2_X1   g498(.A(new_n697), .B(new_n699), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g499(.A(new_n689), .ZN(new_n701));
  INV_X1    g500(.A(new_n538), .ZN(new_n702));
  AOI21_X1  g501(.A(G15gat), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n542), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n701), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n567), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n687), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n631), .A2(new_n664), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT107), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n590), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n693), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n716));
  INV_X1    g515(.A(new_n631), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OR3_X1    g519(.A1(new_n543), .A2(new_n544), .A3(new_n581), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n583), .B1(new_n481), .B2(new_n486), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT35), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n585), .A2(new_n723), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n722), .A2(new_n723), .B1(new_n480), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n720), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n514), .A2(new_n542), .A3(new_n580), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n728), .B2(new_n631), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n663), .B(KEYINPUT108), .Z(new_n731));
  NOR3_X1   g530(.A1(new_n731), .A2(new_n300), .A3(new_n687), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n693), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n734), .A3(new_n735), .ZN(G1328gat));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n733), .B2(new_n391), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n730), .A2(KEYINPUT110), .A3(new_n550), .A4(new_n732), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(G36gat), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n590), .A2(new_n713), .ZN(new_n741));
  NAND2_X1  g540(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n209), .A3(new_n550), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n550), .A2(new_n209), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n714), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n740), .A2(new_n743), .A3(new_n746), .ZN(G1329gat));
  OAI21_X1  g546(.A(new_n719), .B1(new_n582), .B2(new_n589), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n728), .A2(new_n631), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n718), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n748), .A2(new_n750), .A3(new_n704), .A4(new_n732), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n741), .A2(new_n223), .A3(new_n702), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(KEYINPUT112), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n751), .A2(new_n756), .A3(G43gat), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n755), .A2(new_n757), .A3(new_n753), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(G1330gat));
  OAI21_X1  g559(.A(new_n224), .B1(new_n714), .B2(new_n567), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n513), .A2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n733), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT48), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n761), .B(new_n765), .C1(new_n733), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1331gat));
  NOR4_X1   g566(.A1(new_n301), .A2(new_n631), .A3(new_n664), .A4(new_n711), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n728), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n693), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g572(.A1(new_n769), .A2(new_n391), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n770), .A2(G71gat), .A3(new_n704), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n769), .A2(new_n538), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(KEYINPUT113), .ZN(new_n781));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n780), .B2(KEYINPUT113), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n567), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT114), .B(G78gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n301), .A2(new_n663), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n711), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n730), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n771), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n514), .A2(new_n542), .A3(new_n580), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n631), .B(new_n789), .C1(new_n589), .C2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n728), .A2(KEYINPUT51), .A3(new_n631), .A4(new_n789), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n796), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n771), .A2(new_n597), .A3(new_n687), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n793), .A2(new_n597), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NAND4_X1  g603(.A1(new_n748), .A2(new_n750), .A3(new_n550), .A4(new_n791), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n598), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n391), .A2(G92gat), .A3(new_n711), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n800), .A2(new_n801), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n799), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n805), .A2(G92gat), .B1(new_n813), .B2(new_n809), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n808), .A2(new_n812), .B1(new_n811), .B2(new_n814), .ZN(G1337gat));
  AND2_X1   g614(.A1(new_n792), .A2(new_n704), .ZN(new_n816));
  INV_X1    g615(.A(G99gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n538), .A2(G99gat), .A3(new_n711), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT117), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n816), .A2(new_n817), .B1(new_n802), .B2(new_n819), .ZN(G1338gat));
  NAND4_X1  g619(.A1(new_n748), .A2(new_n750), .A3(new_n513), .A4(new_n791), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n567), .A2(G106gat), .A3(new_n711), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n800), .A2(new_n801), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n813), .A2(new_n823), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT118), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n821), .A2(G106gat), .B1(new_n813), .B2(new_n823), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n830), .B(new_n831), .C1(new_n825), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(G1339gat));
  OAI211_X1 g633(.A(new_n279), .B(new_n207), .C1(new_n283), .C2(new_n289), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n266), .A2(new_n270), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n251), .B1(new_n836), .B2(new_n250), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n278), .A2(new_n273), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n205), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n835), .A2(new_n687), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n677), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n682), .B1(new_n685), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n683), .B(new_n846), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n841), .B1(new_n300), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n717), .ZN(new_n852));
  INV_X1    g651(.A(new_n850), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n835), .A2(new_n839), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n631), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n731), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n688), .A2(new_n300), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n585), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n391), .A3(new_n771), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n300), .ZN(new_n862));
  MUX2_X1   g661(.A(G113gat), .B(new_n409), .S(new_n862), .Z(G1340gat));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n711), .ZN(new_n864));
  XOR2_X1   g663(.A(KEYINPUT120), .B(G120gat), .Z(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(G1341gat));
  INV_X1    g665(.A(new_n731), .ZN(new_n867));
  OAI21_X1  g666(.A(G127gat), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n663), .A2(new_n397), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n861), .B2(new_n869), .ZN(G1342gat));
  NAND2_X1  g669(.A1(new_n631), .A2(new_n391), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT121), .Z(new_n872));
  NAND4_X1  g671(.A1(new_n860), .A2(new_n399), .A3(new_n771), .A4(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n861), .B2(new_n717), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  OAI21_X1  g675(.A(new_n513), .B1(new_n856), .B2(new_n858), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT123), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n843), .A2(new_n845), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n683), .A3(new_n846), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n291), .B2(new_n299), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n841), .A3(KEYINPUT122), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n281), .A2(new_n290), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n297), .A2(new_n298), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n883), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(new_n840), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n891), .A3(new_n717), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n663), .B1(new_n892), .B2(new_n855), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n513), .B1(new_n893), .B2(new_n858), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n879), .B1(new_n878), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n855), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n885), .A2(new_n841), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n631), .B1(new_n897), .B2(new_n887), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n886), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n857), .B1(new_n899), .B2(new_n663), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(KEYINPUT123), .A3(KEYINPUT57), .A4(new_n513), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n693), .A2(new_n704), .A3(new_n550), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G141gat), .B1(new_n903), .B2(new_n300), .ZN(new_n904));
  INV_X1    g703(.A(new_n877), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n902), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n419), .A3(new_n301), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT58), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT58), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1344gat));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n901), .A3(new_n687), .A4(new_n902), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n417), .A2(KEYINPUT59), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n913), .A2(KEYINPUT124), .A3(new_n914), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT57), .B1(new_n900), .B2(new_n513), .ZN(new_n919));
  OAI211_X1 g718(.A(KEYINPUT57), .B(new_n513), .C1(new_n856), .C2(new_n858), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n687), .ZN(new_n923));
  OAI21_X1  g722(.A(G148gat), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT59), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n918), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n417), .A3(new_n687), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n903), .B2(new_n867), .ZN(new_n929));
  INV_X1    g728(.A(G155gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n906), .A2(new_n930), .A3(new_n663), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1346gat));
  OAI21_X1  g731(.A(G162gat), .B1(new_n903), .B2(new_n717), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n704), .A2(G162gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n771), .A2(new_n872), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n877), .B2(new_n935), .ZN(G1347gat));
  NOR3_X1   g735(.A1(new_n771), .A2(new_n583), .A3(new_n391), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n859), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n335), .A3(new_n300), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(KEYINPUT125), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n301), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n941), .B2(new_n335), .ZN(G1348gat));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n336), .A3(new_n687), .ZN(new_n943));
  OAI21_X1  g742(.A(G176gat), .B1(new_n938), .B2(new_n711), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  INV_X1    g744(.A(new_n938), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(new_n349), .A3(new_n663), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n342), .B1(new_n946), .B2(new_n731), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  OAI22_X1  g748(.A1(new_n947), .A2(new_n948), .B1(new_n949), .B2(KEYINPUT60), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n938), .B2(new_n717), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT61), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n940), .A2(new_n346), .A3(new_n631), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1351gat));
  NAND3_X1  g755(.A1(new_n693), .A2(new_n550), .A3(new_n542), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n877), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n301), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n894), .A2(new_n878), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n957), .B1(new_n960), .B2(new_n920), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n301), .A2(G197gat), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(new_n961), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n964), .B2(new_n711), .ZN(new_n965));
  NOR4_X1   g764(.A1(new_n877), .A2(new_n957), .A3(G204gat), .A4(new_n711), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n958), .A2(new_n303), .A3(new_n663), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  AOI211_X1 g769(.A(new_n970), .B(new_n303), .C1(new_n961), .C2(new_n663), .ZN(new_n971));
  INV_X1    g770(.A(new_n957), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n663), .B(new_n972), .C1(new_n919), .C2(new_n921), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(KEYINPUT127), .B(new_n969), .C1(new_n971), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(G218gat), .B1(new_n964), .B2(new_n717), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n958), .A2(new_n304), .A3(new_n631), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


