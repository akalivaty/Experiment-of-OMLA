//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT12), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT87), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G104), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(KEYINPUT87), .A3(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(KEYINPUT86), .A3(G104), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n196), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .A4(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n195), .B2(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n195), .A2(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n200), .A2(new_n210), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT88), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n202), .A2(new_n204), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT67), .B(G128), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n205), .B1(G143), .B2(new_n201), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n220), .B(KEYINPUT68), .C1(new_n221), .C2(new_n222), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n206), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n200), .A2(new_n217), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n219), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n226), .A2(new_n206), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n229), .A3(new_n232), .A4(new_n225), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(G137), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n236), .A2(new_n238), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT65), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n242), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n233), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n190), .B1(new_n230), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n229), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT88), .B(new_n218), .C1(new_n248), .C2(new_n227), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT12), .A3(new_n245), .A4(new_n233), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(KEYINPUT89), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G140), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT84), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT74), .B(G953), .Z(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G227), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n253), .B(new_n257), .Z(new_n258));
  AOI22_X1  g072(.A1(new_n212), .A2(new_n213), .B1(new_n195), .B2(G107), .ZN(new_n259));
  OAI21_X1  g073(.A(G101), .B1(new_n259), .B2(KEYINPUT85), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(KEYINPUT85), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT4), .B(new_n217), .C1(new_n265), .C2(new_n260), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n209), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT64), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n209), .A2(new_n271), .A3(KEYINPUT0), .A4(G128), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n245), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT10), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n218), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n248), .A2(new_n227), .A3(KEYINPUT10), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n274), .A2(new_n275), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n190), .C1(new_n230), .C2(new_n246), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n251), .A2(new_n258), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n279), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n258), .A4(new_n251), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n245), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n258), .B1(new_n288), .B2(new_n279), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n258), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n295), .A3(new_n251), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(new_n279), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n258), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G469), .B1(new_n299), .B2(G902), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n189), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT99), .ZN(new_n303));
  INV_X1    g117(.A(G217), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n187), .A2(new_n304), .A3(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n221), .A2(G143), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n203), .A2(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n235), .ZN(new_n310));
  OR2_X1    g124(.A1(KEYINPUT71), .A2(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT71), .A2(G116), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(G122), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n313), .B(new_n192), .C1(new_n314), .C2(G122), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n307), .A2(G134), .A3(new_n308), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n310), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT98), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n311), .A2(KEYINPUT14), .A3(G122), .A4(new_n312), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n319), .A2(G107), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT14), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n313), .B(new_n321), .C1(new_n314), .C2(G122), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n318), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n317), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT97), .B(KEYINPUT13), .Z(new_n327));
  NAND2_X1  g141(.A1(new_n307), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n309), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n328), .A2(G134), .A3(new_n308), .A4(new_n307), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n313), .B1(new_n314), .B2(G122), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n330), .A2(new_n331), .B1(new_n333), .B2(new_n315), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n306), .B1(new_n326), .B2(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n310), .A2(new_n315), .A3(new_n316), .ZN(new_n336));
  INV_X1    g150(.A(new_n325), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n323), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n331), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n315), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n341), .A3(new_n305), .ZN(new_n342));
  AOI21_X1  g156(.A(G902), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G478), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT15), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI211_X1 g161(.A(G902), .B(new_n345), .C1(new_n335), .C2(new_n342), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n303), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n326), .A2(new_n334), .A3(new_n306), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n305), .B1(new_n338), .B2(new_n341), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n293), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n345), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n343), .A2(new_n346), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(KEYINPUT99), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G475), .A2(G902), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT95), .B1(KEYINPUT94), .B2(G143), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(KEYINPUT95), .B2(G143), .ZN(new_n359));
  INV_X1    g173(.A(G237), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n254), .A2(new_n359), .A3(G214), .A4(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(KEYINPUT74), .A2(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT74), .A2(G953), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(G214), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n358), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n239), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT17), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n239), .A3(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G125), .ZN(new_n372));
  INV_X1    g186(.A(G125), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G140), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n374), .A3(KEYINPUT79), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n373), .A2(KEYINPUT79), .A3(G140), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT16), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n377), .A2(new_n201), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n201), .B1(new_n377), .B2(new_n379), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n366), .A2(KEYINPUT17), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n370), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(KEYINPUT18), .A2(G131), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n361), .A2(new_n385), .A3(new_n365), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n375), .A2(new_n376), .A3(G146), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n372), .A2(new_n374), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n201), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n361), .A2(new_n365), .ZN(new_n391));
  INV_X1    g205(.A(new_n385), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT96), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT96), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n394), .B(new_n385), .C1(new_n361), .C2(new_n365), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n386), .B(new_n390), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n195), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n384), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n381), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT19), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n375), .B2(new_n376), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n388), .A2(KEYINPUT19), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n369), .ZN(new_n405));
  OAI221_X1 g219(.A(new_n400), .B1(new_n404), .B2(G146), .C1(new_n405), .C2(new_n366), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n398), .B1(new_n396), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n357), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT20), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n406), .ZN(new_n410));
  INV_X1    g224(.A(new_n398), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n384), .A2(new_n396), .A3(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n357), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n398), .B1(new_n384), .B2(new_n396), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n293), .B1(new_n399), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n409), .A2(new_n416), .B1(G475), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n356), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G214), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(G952), .ZN(new_n422));
  AOI211_X1 g236(.A(G953), .B(new_n422), .C1(G234), .C2(G237), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n293), .B(new_n254), .C1(G234), .C2(G237), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(G898), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(KEYINPUT2), .A2(G113), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT69), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT2), .A2(G113), .ZN(new_n430));
  OR2_X1    g244(.A1(KEYINPUT70), .A2(G119), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT70), .A2(G119), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(G116), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n311), .A2(G119), .A3(new_n312), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n429), .A2(new_n430), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n435), .A2(new_n217), .A3(new_n200), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n433), .A2(KEYINPUT5), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(G113), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(KEYINPUT91), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n437), .A2(new_n438), .A3(new_n442), .A4(G113), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n441), .A2(new_n435), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n444), .B2(new_n248), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT92), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT8), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n270), .A2(new_n272), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n449), .B(G125), .C1(new_n450), .C2(new_n268), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n228), .A2(new_n373), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT93), .B1(new_n273), .B2(new_n373), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G953), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G224), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n445), .A2(new_n448), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n429), .A2(new_n430), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n433), .A2(new_n434), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n435), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n264), .A2(new_n266), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n436), .A2(new_n441), .A3(new_n443), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n447), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n460), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G210), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(G224), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n454), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n467), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n476));
  INV_X1    g290(.A(new_n447), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n477), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n470), .A2(new_n471), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n471), .B1(new_n470), .B2(new_n481), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n421), .B(new_n427), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n302), .A2(new_n420), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT22), .B(G137), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n400), .A2(new_n389), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT23), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n431), .A2(G128), .A3(new_n432), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G128), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n496), .A3(G119), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n492), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n431), .A2(new_n432), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT23), .B1(new_n499), .B2(new_n207), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n498), .A2(new_n500), .A3(G110), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(new_n497), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT24), .B(G110), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(KEYINPUT80), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n498), .ZN(new_n505));
  INV_X1    g319(.A(G110), .ZN(new_n506));
  INV_X1    g320(.A(new_n500), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT80), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n491), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n380), .A2(new_n381), .B1(new_n502), .B2(new_n503), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT78), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(G110), .C1(new_n498), .C2(new_n500), .ZN(new_n514));
  OAI21_X1  g328(.A(G110), .B1(new_n498), .B2(new_n500), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT78), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n490), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n491), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n502), .A2(new_n503), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n508), .B2(new_n509), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n501), .A2(KEYINPUT80), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n512), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n526), .A3(new_n489), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n518), .A2(new_n293), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n518), .A2(new_n527), .A3(new_n293), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n304), .B1(G234), .B2(new_n293), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT77), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT82), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(KEYINPUT82), .A3(new_n536), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n518), .ZN(new_n542));
  INV_X1    g356(.A(new_n527), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT83), .B1(new_n518), .B2(new_n527), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n540), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n237), .A2(KEYINPUT66), .A3(G134), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT66), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n235), .B2(G137), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n237), .A2(G134), .ZN(new_n552));
  OAI211_X1 g366(.A(G131), .B(new_n549), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n241), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n241), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n227), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n242), .A2(G131), .A3(new_n243), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n244), .A2(KEYINPUT65), .A3(new_n241), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n273), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT73), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n227), .A2(new_n563), .A3(new_n555), .A4(new_n557), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(KEYINPUT30), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n227), .A2(new_n241), .A3(new_n553), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n567), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n465), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n465), .B1(new_n245), .B2(new_n273), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n559), .A2(new_n571), .A3(new_n564), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n254), .A2(G210), .A3(new_n360), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT27), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT26), .B(G101), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT75), .B(KEYINPUT31), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n570), .A2(new_n572), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT28), .B1(new_n571), .B2(new_n558), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n567), .A2(new_n562), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n465), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n583), .B2(KEYINPUT28), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n584), .A2(new_n576), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n569), .B1(new_n565), .B2(KEYINPUT30), .ZN(new_n586));
  INV_X1    g400(.A(new_n465), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n572), .B(new_n576), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  OR2_X1    g402(.A1(KEYINPUT75), .A2(KEYINPUT31), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(G472), .A2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT32), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n572), .B1(new_n586), .B2(new_n587), .ZN(new_n598));
  INV_X1    g412(.A(new_n576), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(KEYINPUT76), .A3(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT29), .B1(new_n584), .B2(new_n576), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT28), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n565), .A2(new_n465), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(new_n572), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n580), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n576), .A2(KEYINPUT29), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n548), .B1(new_n597), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n486), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n591), .A2(new_n293), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(G472), .B1(new_n591), .B2(new_n592), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n534), .A2(KEYINPUT82), .A3(new_n536), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT82), .B1(new_n534), .B2(new_n536), .ZN(new_n620));
  INV_X1    g434(.A(new_n547), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n622), .A3(new_n301), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT100), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n618), .A2(new_n622), .A3(new_n625), .A4(new_n301), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n418), .A2(G475), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n415), .B1(new_n414), .B2(new_n357), .ZN(new_n628));
  INV_X1    g442(.A(new_n357), .ZN(new_n629));
  AOI211_X1 g443(.A(KEYINPUT20), .B(new_n629), .C1(new_n412), .C2(new_n413), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n627), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT33), .B1(new_n350), .B2(new_n351), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n335), .A2(new_n342), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(G478), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n344), .A2(new_n293), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n343), .B2(new_n344), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(KEYINPUT101), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n485), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n624), .A2(new_n626), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT102), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NOR3_X1   g460(.A1(new_n485), .A2(new_n631), .A3(new_n356), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n624), .A2(new_n626), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NAND2_X1  g464(.A1(new_n523), .A2(new_n526), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n490), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n541), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n539), .A2(new_n540), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n618), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n486), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  XOR2_X1   g473(.A(KEYINPUT103), .B(G900), .Z(new_n660));
  AOI21_X1  g474(.A(new_n423), .B1(new_n424), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n419), .A2(new_n355), .A3(new_n349), .A4(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n301), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n666));
  INV_X1    g480(.A(new_n596), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n613), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n421), .ZN(new_n669));
  INV_X1    g483(.A(new_n471), .ZN(new_n670));
  INV_X1    g484(.A(new_n481), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n445), .A2(new_n448), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n455), .A2(new_n459), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n461), .A2(new_n468), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n293), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n670), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n669), .B1(new_n677), .B2(new_n482), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n665), .A2(new_n668), .A3(new_n678), .A4(new_n655), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n482), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n655), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n356), .A2(new_n419), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n421), .A2(new_n683), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n661), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n301), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n598), .A2(new_n576), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n607), .A2(new_n572), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n691), .B(new_n293), .C1(new_n576), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G472), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n667), .B2(new_n666), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n686), .A2(new_n689), .A3(new_n690), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT105), .B(G143), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G45));
  NAND3_X1  g512(.A1(new_n631), .A2(new_n638), .A3(new_n662), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n189), .B(new_n699), .C1(new_n294), .C2(new_n300), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n668), .A2(new_n700), .A3(new_n678), .A4(new_n655), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NAND2_X1  g516(.A1(new_n294), .A2(new_n188), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n291), .A2(new_n293), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n292), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n289), .B1(new_n282), .B2(KEYINPUT90), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n707), .B2(new_n286), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n703), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n668), .A2(new_n642), .A3(new_n710), .A4(new_n622), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND4_X1  g527(.A1(new_n668), .A2(new_n710), .A3(new_n647), .A4(new_n622), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AOI21_X1  g529(.A(new_n189), .B1(new_n708), .B2(new_n292), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n708), .B2(KEYINPUT106), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n705), .B(G902), .C1(new_n707), .C2(new_n286), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n678), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n704), .A2(new_n705), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(G469), .A3(new_n709), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(KEYINPUT107), .A3(new_n678), .A4(new_n716), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(G472), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n605), .B2(new_n611), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n594), .B2(new_n596), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n420), .A2(new_n426), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n728), .A2(new_n684), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NAND2_X1  g547(.A1(new_n548), .A2(KEYINPUT109), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n539), .A2(new_n735), .A3(new_n540), .A4(new_n547), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n617), .A2(G472), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT108), .B1(new_n608), .B2(new_n580), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n599), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n608), .A2(KEYINPUT108), .A3(new_n580), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n579), .A2(new_n590), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n592), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n485), .A2(new_n419), .A3(new_n356), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n737), .A2(new_n710), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  INV_X1    g562(.A(new_n699), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n655), .A2(new_n738), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n725), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n725), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  NOR3_X1   g571(.A1(new_n483), .A2(new_n669), .A3(new_n484), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n749), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n302), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n737), .A3(new_n668), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n301), .A2(new_n758), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n728), .A2(new_n762), .A3(new_n548), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n761), .A2(KEYINPUT42), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  XOR2_X1   g580(.A(new_n663), .B(KEYINPUT111), .Z(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  OAI21_X1  g583(.A(G469), .B1(new_n299), .B2(KEYINPUT45), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT112), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n770), .A2(KEYINPUT112), .B1(KEYINPUT45), .B2(new_n299), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(G469), .A2(G902), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT46), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n292), .B2(new_n708), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n774), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n189), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n687), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n684), .A2(new_n618), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n419), .A2(new_n638), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT43), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n631), .B2(KEYINPUT113), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n783), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n780), .A2(new_n758), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NOR2_X1   g607(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n778), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n778), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n668), .A2(new_n622), .A3(new_n759), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NAND4_X1  g615(.A1(new_n737), .A2(new_n188), .A3(new_n421), .A4(new_n783), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n723), .A2(new_n294), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n803), .A2(KEYINPUT116), .B1(KEYINPUT49), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n695), .B(new_n683), .C1(new_n802), .C2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n805), .B(new_n807), .C1(KEYINPUT49), .C2(new_n804), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n678), .A2(new_n662), .A3(new_n685), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n655), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n301), .A3(new_n695), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n679), .A2(new_n701), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n754), .B1(new_n725), .B2(new_n751), .ZN(new_n813));
  AOI211_X1 g627(.A(KEYINPUT110), .B(new_n750), .C1(new_n721), .C2(new_n724), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n812), .B(KEYINPUT52), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n747), .A2(new_n711), .A3(new_n714), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n667), .A2(new_n666), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n729), .B(new_n655), .C1(new_n823), .C2(new_n727), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n721), .B2(new_n724), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n614), .B(new_n710), .C1(new_n642), .C2(new_n647), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n732), .A2(new_n827), .A3(new_n747), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n347), .A2(new_n348), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n631), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n832), .A2(KEYINPUT118), .B1(new_n631), .B2(new_n638), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n485), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n624), .A2(new_n626), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n486), .B1(new_n614), .B2(new_n656), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n419), .A2(new_n831), .A3(new_n662), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n668), .A2(new_n655), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n750), .ZN(new_n841));
  INV_X1    g655(.A(new_n762), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n838), .A2(new_n765), .A3(new_n768), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n830), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n817), .A2(KEYINPUT119), .A3(new_n818), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n821), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n819), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n763), .A2(new_n764), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n843), .A2(new_n852), .A3(new_n853), .A4(new_n768), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n732), .A2(KEYINPUT53), .A3(new_n747), .A4(new_n828), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n836), .A2(new_n837), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(new_n756), .B2(new_n812), .ZN(new_n858));
  INV_X1    g672(.A(new_n818), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n819), .A2(KEYINPUT120), .A3(new_n857), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n846), .A2(new_n845), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT119), .B1(new_n817), .B2(new_n818), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n849), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n864), .A2(new_n867), .A3(KEYINPUT121), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n851), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n847), .A2(new_n849), .B1(new_n862), .B2(new_n863), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n871), .B2(new_n868), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n786), .A2(new_n423), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT122), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n737), .A2(new_n745), .ZN(new_n876));
  INV_X1    g690(.A(new_n710), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n683), .A3(new_n421), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT50), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n875), .A2(new_n710), .A3(new_n758), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n745), .A2(new_n655), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n710), .A2(new_n758), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n622), .A2(new_n423), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n695), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n631), .A2(new_n638), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n881), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n875), .A2(new_n876), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n758), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n796), .A2(new_n798), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n723), .A2(new_n189), .A3(new_n294), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n873), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n798), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n795), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n758), .A3(new_n892), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n885), .A2(new_n890), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(KEYINPUT51), .A3(new_n881), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n892), .A2(new_n725), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n640), .A2(new_n641), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n422), .B(G953), .C1(new_n888), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n728), .B1(new_n734), .B2(new_n736), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n882), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(KEYINPUT48), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(KEYINPUT48), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n897), .A2(new_n902), .A3(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n870), .A2(new_n872), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n808), .B1(new_n913), .B2(new_n914), .ZN(G75));
  AOI21_X1  g729(.A(new_n293), .B1(new_n864), .B2(new_n867), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(G210), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n480), .A2(new_n478), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n474), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n671), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n917), .B2(new_n918), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n254), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  NOR4_X1   g740(.A1(new_n871), .A2(KEYINPUT123), .A3(new_n293), .A4(new_n773), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n928));
  INV_X1    g742(.A(new_n773), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n916), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n774), .B(KEYINPUT57), .Z(new_n932));
  AND3_X1   g746(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n868), .B1(new_n864), .B2(new_n867), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n291), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n925), .B1(new_n931), .B2(new_n936), .ZN(G54));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n916), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n414), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n939), .A2(KEYINPUT124), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n916), .A2(new_n414), .A3(new_n938), .ZN(new_n943));
  INV_X1    g757(.A(new_n925), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(G60));
  AND2_X1   g760(.A1(new_n632), .A2(new_n634), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n636), .B(KEYINPUT59), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n933), .B2(new_n934), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n944), .ZN(new_n951));
  INV_X1    g765(.A(new_n948), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n870), .B2(new_n872), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n947), .B2(new_n953), .ZN(G63));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n925), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT60), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n864), .B2(new_n867), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n545), .A2(new_n546), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n958), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n653), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n871), .A2(new_n965), .A3(new_n960), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n957), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n962), .B1(new_n871), .B2(new_n960), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n961), .A2(new_n653), .ZN(new_n969));
  INV_X1    g783(.A(new_n957), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n958), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n967), .A2(new_n971), .ZN(G66));
  NAND3_X1  g786(.A1(new_n826), .A2(new_n829), .A3(new_n838), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n254), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n425), .B2(new_n472), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(G898), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n919), .B1(new_n977), .B2(new_n255), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n976), .B(new_n978), .Z(G69));
  NAND2_X1  g793(.A1(new_n833), .A2(new_n834), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n758), .B1(new_n980), .B2(KEYINPUT126), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(KEYINPUT126), .B2(new_n980), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n614), .A3(new_n301), .A4(new_n687), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n792), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n756), .A2(new_n679), .A3(new_n701), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n696), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n985), .A2(new_n988), .A3(new_n696), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n984), .A2(new_n987), .A3(new_n800), .A4(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n990), .A2(new_n254), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n586), .B(new_n404), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n780), .A2(new_n678), .A3(new_n685), .A4(new_n907), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n993), .A2(new_n765), .A3(new_n768), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n994), .A2(new_n792), .A3(new_n800), .A4(new_n985), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n255), .ZN(new_n996));
  INV_X1    g810(.A(G900), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n992), .B1(new_n997), .B2(new_n254), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n991), .A2(new_n992), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n255), .B1(new_n256), .B2(new_n997), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1002), .ZN(new_n1004));
  OAI221_X1 g818(.A(new_n1004), .B1(new_n996), .B2(new_n998), .C1(new_n991), .C2(new_n992), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n995), .B2(new_n973), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n570), .A2(new_n572), .A3(new_n599), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n925), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n602), .A2(new_n603), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n588), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n848), .A2(new_n850), .A3(new_n1008), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1008), .B1(new_n990), .B2(new_n973), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n576), .A3(new_n598), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(G57));
endmodule


