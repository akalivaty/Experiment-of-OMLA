//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(new_n211), .B2(KEYINPUT66), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n207), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G13), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G250), .B1(G257), .B2(G264), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n217), .A2(new_n218), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n219), .B(new_n228), .C1(new_n231), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT67), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G223), .A3(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n252), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(new_n257), .B2(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(new_n264), .ZN(new_n268));
  INV_X1    g0068(.A(G226), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G179), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n203), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n230), .A2(G33), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n274), .B1(new_n275), .B2(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT69), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(new_n282), .B1(G1), .B2(G13), .ZN(new_n283));
  NAND4_X1  g0083(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n280), .A2(new_n285), .B1(new_n202), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(new_n263), .B2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n270), .B1(new_n258), .B2(new_n261), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(G169), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n288), .A2(KEYINPUT9), .A3(new_n290), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n296), .B(new_n297), .C1(new_n292), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(G190), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT10), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n296), .A2(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n272), .A2(G200), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n300), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n294), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n278), .B(KEYINPUT70), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n277), .ZN(new_n309));
  XOR2_X1   g0109(.A(KEYINPUT15), .B(G87), .Z(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n311), .A2(new_n279), .B1(new_n230), .B2(new_n256), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n285), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n286), .A2(G77), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n289), .B2(G77), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n252), .ZN(new_n320));
  INV_X1    g0120(.A(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G232), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n325), .A2(new_n326), .A3(G1698), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n317), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n268), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n266), .B1(new_n329), .B2(G244), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n316), .B1(G190), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n313), .A2(new_n315), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n307), .A2(KEYINPUT71), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n252), .A2(G226), .A3(new_n253), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G97), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n317), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n266), .B1(new_n329), .B2(G238), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G200), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n289), .A2(G68), .ZN(new_n355));
  INV_X1    g0155(.A(G68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n287), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n279), .A2(new_n256), .B1(new_n230), .B2(G68), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(KEYINPUT72), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n277), .B2(new_n202), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n276), .A2(KEYINPUT73), .A3(G50), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(new_n362), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n285), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT11), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n366), .A2(new_n369), .A3(new_n285), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n359), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n350), .A2(G190), .A3(new_n352), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n354), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT74), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n354), .A2(new_n372), .A3(KEYINPUT74), .A4(new_n371), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n353), .B2(G169), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n353), .A2(new_n338), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n353), .A2(new_n378), .A3(G169), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n278), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n287), .ZN(new_n386));
  INV_X1    g0186(.A(new_n289), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n385), .ZN(new_n388));
  INV_X1    g0188(.A(new_n285), .ZN(new_n389));
  INV_X1    g0189(.A(G58), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n356), .ZN(new_n391));
  OAI21_X1  g0191(.A(G20), .B1(new_n391), .B2(new_n201), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n276), .A2(G159), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n323), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT7), .B(new_n230), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n325), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n230), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n252), .B2(G20), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n394), .B1(new_n403), .B2(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n389), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(new_n394), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT76), .B1(new_n321), .B2(KEYINPUT3), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n323), .A3(G33), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n410), .A3(new_n322), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n401), .A2(G20), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n356), .B1(new_n413), .B2(new_n402), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT77), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n325), .A2(new_n230), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n401), .B1(new_n411), .B2(new_n412), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n418), .A2(KEYINPUT77), .A3(new_n356), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n406), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n388), .B1(new_n405), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n322), .A2(new_n324), .A3(G223), .A4(new_n253), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n252), .A2(KEYINPUT78), .A3(G223), .A4(new_n253), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n252), .A2(G226), .A3(G1698), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n317), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n267), .B1(new_n268), .B2(new_n326), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n336), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n338), .B(new_n431), .C1(new_n429), .C2(new_n317), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n421), .A2(new_n422), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n422), .B1(new_n421), .B2(new_n435), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n298), .B1(new_n430), .B2(new_n432), .ZN(new_n441));
  INV_X1    g0241(.A(G190), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n442), .B(new_n431), .C1(new_n429), .C2(new_n317), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n421), .A2(new_n440), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n440), .B1(new_n421), .B2(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n342), .A2(new_n384), .A3(new_n439), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT71), .B1(new_n307), .B2(new_n341), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(G20), .B1(G33), .B2(G283), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n321), .A2(G97), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n453), .A2(new_n454), .B1(G20), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n285), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n285), .A2(KEYINPUT20), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n263), .A2(G33), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n286), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(G116), .A3(new_n284), .A4(new_n283), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n287), .A2(new_n455), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(G303), .B1(new_n395), .B2(new_n396), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n322), .A2(new_n324), .A3(G257), .A4(new_n253), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n322), .A2(new_n324), .A3(G264), .A4(G1698), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n317), .ZN(new_n473));
  INV_X1    g0273(.A(G41), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n263), .B(G45), .C1(new_n474), .C2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G41), .ZN(new_n477));
  OAI211_X1 g0277(.A(G270), .B(new_n260), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n263), .A2(G45), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(G41), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(G274), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n336), .B1(new_n473), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT21), .B1(new_n468), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n478), .A2(new_n483), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n317), .B2(new_n472), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n485), .A2(KEYINPUT21), .B1(new_n489), .B2(G179), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n466), .B1(new_n459), .B2(new_n460), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n489), .A2(new_n493), .A3(new_n336), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n473), .A2(new_n484), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n338), .ZN(new_n496));
  OAI211_X1 g0296(.A(KEYINPUT80), .B(new_n468), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n486), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n287), .A2(new_n319), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n463), .A2(new_n284), .A3(new_n283), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(G107), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(KEYINPUT81), .A2(G87), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n322), .A2(new_n324), .A3(new_n503), .A4(new_n230), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n252), .A2(KEYINPUT22), .A3(new_n230), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G20), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n230), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n319), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n506), .A2(new_n507), .A3(new_n513), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(KEYINPUT24), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n285), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT24), .B1(new_n515), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n502), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n322), .A2(new_n324), .A3(G250), .A4(new_n253), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n322), .A2(new_n324), .A3(G257), .A4(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n475), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n317), .B1(new_n526), .B2(new_n481), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n317), .A2(new_n525), .B1(new_n527), .B2(G264), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n483), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(G179), .ZN(new_n530));
  AOI21_X1  g0330(.A(G169), .B1(new_n528), .B2(new_n483), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n521), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n498), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n298), .B1(new_n528), .B2(new_n483), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n317), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n527), .A2(G264), .ZN(new_n537));
  AND4_X1   g0337(.A1(G190), .A2(new_n536), .A3(new_n537), .A4(new_n483), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n539), .B(new_n502), .C1(new_n520), .C2(new_n519), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n495), .A2(G200), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n473), .A2(new_n484), .A3(G190), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n491), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n322), .A2(new_n324), .A3(G238), .A4(new_n253), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n322), .A2(new_n324), .A3(G244), .A4(G1698), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n508), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n317), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n479), .A2(G250), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n317), .A2(new_n548), .B1(new_n265), .B2(new_n479), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n230), .B1(new_n345), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G87), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n319), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n322), .A2(new_n324), .A3(new_n230), .A4(G68), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n553), .B1(new_n279), .B2(new_n556), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n285), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n463), .A2(G87), .A3(new_n284), .A4(new_n283), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n311), .A2(new_n287), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n549), .B1(new_n546), .B2(new_n317), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n552), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n338), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n463), .A2(new_n310), .A3(new_n284), .A4(new_n283), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n571), .C1(G169), .C2(new_n566), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n543), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n556), .A2(new_n319), .A3(KEYINPUT6), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n319), .A2(KEYINPUT79), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G107), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n574), .A2(new_n576), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n574), .A2(new_n576), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(G20), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n276), .A2(G77), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n418), .C2(new_n319), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n285), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n501), .A2(G97), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n286), .A2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G257), .B(new_n260), .C1(new_n475), .C2(new_n477), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n483), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n322), .A2(new_n324), .A3(G244), .A4(new_n253), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n597));
  NAND2_X1  g0397(.A1(G33), .A2(G283), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n593), .B1(new_n600), .B2(new_n317), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n336), .ZN(new_n603));
  AOI211_X1 g0403(.A(G179), .B(new_n593), .C1(new_n600), .C2(new_n317), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n591), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n589), .B1(new_n285), .B2(new_n584), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(G190), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n298), .C2(new_n601), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n540), .A2(new_n573), .A3(new_n606), .A4(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n452), .A2(new_n534), .A3(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n340), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n383), .B1(new_n612), .B2(new_n373), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n439), .B1(new_n613), .B2(new_n447), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n302), .A2(new_n306), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n294), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n572), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n601), .A2(G169), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n607), .A2(new_n618), .A3(new_n604), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n568), .A2(new_n572), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n617), .B1(new_n621), .B2(KEYINPUT26), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT83), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n551), .A2(new_n623), .A3(G200), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT83), .B1(new_n566), .B2(new_n298), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(new_n567), .A4(new_n565), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n572), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n619), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n495), .A2(KEYINPUT21), .A3(G169), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n489), .A2(G179), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n491), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT84), .B1(new_n633), .B2(new_n486), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n495), .A2(G169), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n493), .B1(new_n635), .B2(new_n491), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT84), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(new_n491), .C2(new_n490), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n533), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n628), .A2(new_n540), .A3(new_n606), .A4(new_n609), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n622), .B(new_n630), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n616), .B1(new_n452), .B2(new_n642), .ZN(G369));
  NOR2_X1   g0443(.A1(new_n220), .A2(G20), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n263), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n491), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n543), .B1(new_n498), .B2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n634), .A2(new_n638), .A3(new_n652), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n498), .B2(new_n650), .ZN(new_n657));
  INV_X1    g0457(.A(new_n533), .ZN(new_n658));
  INV_X1    g0458(.A(new_n540), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n521), .A2(new_n650), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(KEYINPUT85), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n533), .A2(new_n650), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(KEYINPUT86), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n221), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n557), .A2(G116), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G1), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n234), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n669), .B2(new_n673), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT28), .Z(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n628), .A2(new_n606), .A3(new_n609), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n534), .A3(new_n540), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT26), .B1(new_n606), .B2(new_n627), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n619), .A2(new_n620), .A3(new_n629), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n572), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI211_X1 g0484(.A(new_n678), .B(new_n650), .C1(new_n680), .C2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT29), .B1(new_n641), .B2(new_n651), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT88), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n650), .B1(new_n680), .B2(new_n684), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT88), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G330), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n489), .A2(new_n528), .A3(G179), .A4(new_n566), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n602), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n489), .A2(G179), .A3(new_n566), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n529), .A3(new_n602), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n528), .A2(new_n566), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n496), .A3(KEYINPUT30), .A4(new_n601), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT87), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n696), .A2(new_n698), .A3(new_n700), .A4(KEYINPUT87), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n650), .A3(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n534), .A2(new_n610), .A3(new_n650), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n693), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n692), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n677), .B1(new_n713), .B2(G1), .ZN(G364));
  AOI21_X1  g0514(.A(new_n263), .B1(new_n644), .B2(G45), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n671), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n655), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT89), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n229), .B1(G20), .B2(new_n336), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n247), .A2(G45), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n221), .A2(new_n252), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(G45), .C2(new_n233), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n221), .A2(new_n325), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n729), .A2(G355), .B1(new_n455), .B2(new_n221), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n725), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n230), .A2(G190), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(G179), .A3(new_n298), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT91), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n733), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n738), .A2(G283), .B1(G329), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n230), .A2(new_n442), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n338), .A2(new_n298), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n252), .B1(new_n746), .B2(G326), .ZN(new_n747));
  INV_X1    g0547(.A(new_n743), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n298), .A3(G179), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n338), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n732), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n749), .A2(G303), .B1(G311), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n744), .A2(new_n732), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT33), .B(G317), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n743), .A2(new_n750), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(new_n756), .B1(new_n758), .B2(G322), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n742), .A2(new_n747), .A3(new_n753), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(G20), .B1(new_n740), .B2(new_n442), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n738), .A2(G107), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n325), .B1(new_n746), .B2(G50), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n749), .A2(G87), .B1(G77), .B2(new_n752), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G58), .A2(new_n758), .B1(new_n755), .B2(G68), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n741), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT32), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n762), .C2(new_n556), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n760), .A2(new_n764), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n731), .B1(new_n775), .B2(new_n723), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n716), .B1(new_n722), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n716), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n717), .A2(new_n693), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n779), .B2(new_n656), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  NOR2_X1   g0583(.A1(new_n340), .A2(new_n650), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n316), .A2(new_n650), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n335), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(new_n786), .B2(new_n340), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n642), .B2(new_n650), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n641), .A2(new_n651), .A3(new_n787), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n711), .A2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT96), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT96), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n778), .B1(new_n711), .B2(new_n791), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n723), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n738), .A2(G68), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n325), .B1(new_n749), .B2(G50), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n770), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G58), .B2(new_n761), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n802), .A2(KEYINPUT94), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n746), .A2(G137), .B1(new_n752), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(G143), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n805), .B2(new_n757), .C1(new_n275), .C2(new_n754), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT34), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n802), .B2(KEYINPUT94), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n738), .A2(G87), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n770), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT93), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n746), .A2(G303), .B1(new_n752), .B2(G116), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n814), .B2(new_n754), .C1(new_n763), .C2(new_n757), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n252), .B(new_n815), .C1(G107), .C2(new_n749), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n556), .B2(new_n762), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n803), .A2(new_n808), .B1(new_n812), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n797), .B1(new_n818), .B2(KEYINPUT95), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(KEYINPUT95), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n723), .A2(new_n718), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n716), .B1(new_n256), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(new_n720), .C2(new_n787), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n796), .A2(new_n823), .ZN(G384));
  OAI21_X1  g0624(.A(G77), .B1(new_n390), .B2(new_n356), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n233), .A2(new_n825), .B1(G50), .B2(new_n356), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(G1), .A3(new_n220), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n580), .A2(new_n581), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(KEYINPUT35), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(G116), .A3(new_n231), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(KEYINPUT35), .B2(new_n830), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n828), .B1(new_n833), .B2(KEYINPUT36), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(KEYINPUT36), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n644), .A2(new_n263), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n405), .A2(new_n420), .ZN(new_n837));
  INV_X1    g0637(.A(new_n388), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n837), .A2(new_n838), .A3(new_n444), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT7), .B1(new_n325), .B2(new_n230), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n398), .B2(new_n397), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n356), .B1(new_n841), .B2(new_n400), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n406), .B1(new_n842), .B2(new_n394), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n405), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(new_n838), .B1(new_n435), .B2(new_n648), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT37), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n837), .A2(new_n838), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n435), .A2(new_n648), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n421), .A2(new_n444), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT98), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n846), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n846), .B2(new_n852), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n438), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n436), .B1(new_n445), .B2(new_n446), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n648), .B1(new_n844), .B2(new_n838), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n846), .A2(new_n852), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT98), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n846), .A2(new_n852), .A3(new_n853), .ZN(new_n864));
  AND4_X1   g0664(.A1(KEYINPUT38), .A2(new_n863), .A3(new_n860), .A4(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT39), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(new_n648), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n847), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n448), .B2(new_n439), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n849), .A2(new_n851), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(new_n850), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n863), .A2(new_n860), .A3(KEYINPUT38), .A4(new_n864), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n381), .A2(new_n382), .ZN(new_n878));
  INV_X1    g0678(.A(new_n371), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n650), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT99), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n863), .A2(new_n860), .A3(new_n864), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n867), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n874), .ZN(new_n887));
  INV_X1    g0687(.A(new_n784), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n790), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n371), .A2(new_n651), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n375), .A2(new_n376), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n880), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n373), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n383), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n887), .B(new_n890), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n439), .B2(new_n868), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n687), .A2(new_n451), .A3(new_n691), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n616), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n899), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n705), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n492), .A2(new_n497), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n904), .A2(new_n533), .A3(new_n636), .ZN(new_n905));
  AND4_X1   g0705(.A1(new_n540), .A2(new_n573), .A3(new_n606), .A4(new_n609), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n651), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n903), .B1(new_n907), .B2(KEYINPUT31), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n705), .A2(new_n707), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n787), .B1(new_n894), .B2(new_n896), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n887), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n873), .A2(new_n874), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n916), .B2(new_n913), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(G330), .ZN(new_n918));
  INV_X1    g0718(.A(new_n909), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n693), .B1(new_n708), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n451), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n452), .A2(new_n910), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n918), .A2(new_n921), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n836), .B1(new_n902), .B2(new_n923), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n924), .A2(KEYINPUT100), .B1(new_n902), .B2(new_n923), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(KEYINPUT100), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n835), .B1(new_n925), .B2(new_n926), .ZN(G367));
  NOR2_X1   g0727(.A1(new_n498), .A2(new_n650), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n665), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n609), .B(new_n606), .C1(new_n607), .C2(new_n651), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT42), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n619), .A2(new_n650), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT101), .Z(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(new_n533), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n606), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT102), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT102), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n940), .A3(new_n606), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n651), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT43), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n651), .A2(new_n565), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n628), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n572), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n933), .A2(new_n942), .A3(new_n943), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n943), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n939), .A2(new_n651), .A3(new_n941), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n932), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n656), .A2(new_n663), .A3(new_n664), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n936), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n949), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n956), .B1(new_n949), .B2(new_n953), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n715), .B(KEYINPUT103), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n929), .A2(new_n667), .A3(new_n935), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT45), .Z(new_n963));
  AOI21_X1  g0763(.A(new_n935), .B1(new_n929), .B2(new_n667), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT44), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n955), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n657), .B(new_n665), .Z(new_n967));
  AOI21_X1  g0767(.A(new_n712), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n670), .B(KEYINPUT41), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n961), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n948), .A2(new_n721), .ZN(new_n972));
  INV_X1    g0772(.A(new_n221), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n724), .B1(new_n973), .B2(new_n311), .ZN(new_n974));
  INV_X1    g0774(.A(new_n727), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n242), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n778), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  INV_X1    g0778(.A(new_n749), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n455), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n749), .A2(KEYINPUT46), .A3(G116), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n252), .B1(new_n746), .B2(G311), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G107), .B2(new_n761), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G303), .A2(new_n758), .B1(new_n752), .B2(G283), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n763), .B2(new_n754), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n738), .B2(G97), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n984), .B(new_n987), .C1(new_n988), .C2(new_n770), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n738), .A2(G77), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n252), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT104), .Z(new_n992));
  AOI22_X1  g0792(.A1(new_n749), .A2(G58), .B1(G150), .B2(new_n758), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n771), .B2(new_n754), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n745), .A2(new_n805), .B1(new_n751), .B2(new_n202), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n761), .A2(G68), .ZN(new_n997));
  INV_X1    g0797(.A(G137), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n997), .C1(new_n998), .C2(new_n770), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n989), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT47), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n797), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n977), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n959), .A2(new_n971), .B1(new_n972), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT105), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(KEYINPUT105), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(G387));
  NAND2_X1  g0810(.A1(new_n713), .A2(new_n967), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n671), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n713), .B2(new_n967), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n721), .B1(new_n663), .B2(new_n664), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n672), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n729), .A2(new_n1016), .B1(new_n319), .B2(new_n221), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT106), .Z(new_n1018));
  NOR2_X1   g0818(.A1(new_n308), .A2(G50), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n1016), .C1(G68), .C2(G77), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n975), .B1(new_n239), .B2(G45), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n778), .B1(new_n1026), .B2(new_n725), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n979), .A2(new_n256), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G68), .B2(new_n752), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n202), .B2(new_n757), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G97), .B2(new_n738), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n746), .A2(G159), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT107), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n252), .B1(new_n278), .B2(new_n754), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n762), .A2(new_n311), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n1033), .C2(new_n1032), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1031), .B(new_n1036), .C1(new_n275), .C2(new_n770), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n746), .A2(G322), .B1(new_n752), .B2(G303), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n810), .B2(new_n754), .C1(new_n988), .C2(new_n757), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT48), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n814), .B2(new_n762), .C1(new_n763), .C2(new_n979), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT49), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n741), .A2(G326), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n325), .B(new_n1043), .C1(new_n737), .C2(new_n455), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1037), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1027), .B1(new_n1045), .B2(new_n723), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n967), .A2(new_n960), .B1(new_n1015), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1014), .A2(new_n1047), .ZN(G393));
  AOI21_X1  g0848(.A(new_n955), .B1(new_n963), .B2(new_n965), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(KEYINPUT108), .A3(new_n966), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n966), .A2(KEYINPUT108), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n1049), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n961), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n755), .A2(G303), .B1(new_n752), .B2(G294), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n745), .A2(new_n988), .B1(new_n757), .B2(new_n810), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT111), .Z(new_n1057));
  OAI221_X1 g0857(.A(new_n1055), .B1(new_n455), .B2(new_n762), .C1(new_n1057), .C2(KEYINPUT52), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n741), .A2(G322), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n252), .B1(new_n749), .B2(G283), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n765), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT112), .Z(new_n1062));
  AOI211_X1 g0862(.A(new_n1058), .B(new_n1062), .C1(KEYINPUT52), .C2(new_n1057), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n252), .B1(new_n979), .B2(new_n356), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G50), .B2(new_n755), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n809), .B(new_n1065), .C1(new_n256), .C2(new_n762), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n745), .A2(new_n275), .B1(new_n757), .B2(new_n771), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1068));
  XNOR2_X1  g0868(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n770), .A2(new_n805), .B1(new_n308), .B2(new_n751), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1066), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT110), .Z(new_n1072));
  OAI21_X1  g0872(.A(new_n723), .B1(new_n1063), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n936), .A2(new_n721), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n725), .B1(G97), .B2(new_n221), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n975), .A2(new_n250), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n716), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1073), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1054), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1051), .A2(new_n1011), .A3(new_n1053), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n671), .B1(new_n966), .B2(new_n1012), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(new_n709), .ZN(new_n1085));
  OAI211_X1 g0885(.A(G330), .B(new_n787), .C1(new_n908), .C2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n894), .A2(new_n896), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n896), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n891), .B1(new_n377), .B2(new_n383), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n788), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n920), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(G330), .B1(new_n908), .B2(new_n909), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1087), .B1(new_n1094), .B2(new_n788), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n786), .A2(new_n340), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n905), .A2(new_n640), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n651), .B(new_n1096), .C1(new_n1097), .C2(new_n683), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n888), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n710), .B2(new_n1091), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1093), .A2(new_n890), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n900), .A2(new_n616), .A3(new_n921), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT114), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1095), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1087), .A2(new_n1086), .B1(new_n920), .B2(new_n1091), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n889), .B2(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n900), .A2(new_n616), .A3(new_n921), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT114), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n883), .B1(new_n889), .B2(new_n1087), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n866), .A2(new_n876), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1099), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n915), .B(new_n883), .C1(new_n1087), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n710), .A2(new_n1091), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT113), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT113), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1112), .A2(new_n1118), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1092), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n671), .B1(new_n1110), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT115), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1116), .A2(KEYINPUT113), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1128));
  AND4_X1   g0928(.A1(KEYINPUT115), .A2(new_n1126), .A3(new_n1128), .A4(new_n1119), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n877), .A2(new_n719), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n821), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n778), .B1(new_n385), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g0933(.A(KEYINPUT54), .B(G143), .Z(new_n1134));
  AOI22_X1  g0934(.A1(new_n755), .A2(G137), .B1(new_n752), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n762), .B2(new_n771), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT116), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n252), .B1(new_n757), .B2(new_n800), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G128), .B2(new_n746), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n749), .A2(G150), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT53), .Z(new_n1141));
  AOI22_X1  g0941(.A1(new_n738), .A2(G50), .B1(G125), .B2(new_n741), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n798), .B(new_n325), .C1(new_n555), .C2(new_n979), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G294), .B2(new_n741), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n762), .A2(new_n256), .B1(new_n455), .B2(new_n757), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n745), .A2(new_n814), .B1(new_n751), .B2(new_n556), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G107), .B2(new_n755), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT117), .Z(new_n1150));
  NAND3_X1  g0950(.A1(new_n1145), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1143), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1133), .B1(new_n1153), .B2(new_n723), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1125), .A2(new_n960), .B1(new_n1131), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1130), .A2(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(new_n294), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n615), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT55), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n307), .A2(KEYINPUT55), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n291), .A2(new_n868), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(new_n1163), .A3(new_n1161), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n918), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT120), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1166), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(KEYINPUT120), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n917), .A3(G330), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1171), .A2(KEYINPUT121), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n899), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n897), .B1(new_n439), .B2(new_n868), .C1(new_n877), .C2(new_n883), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1171), .A2(new_n1183), .A3(KEYINPUT121), .A4(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n960), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n738), .A2(G58), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n325), .A2(new_n474), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n311), .A2(new_n751), .B1(new_n319), .B2(new_n757), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n745), .A2(new_n455), .B1(new_n754), .B2(new_n556), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1028), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n741), .A2(G283), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1187), .A2(new_n1191), .A3(new_n997), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT58), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1188), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G128), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n757), .A2(new_n1198), .B1(new_n751), .B2(new_n998), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G125), .B2(new_n746), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n749), .A2(new_n1134), .B1(G132), .B2(new_n755), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n275), .C2(new_n762), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n738), .A2(G159), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n741), .C2(G124), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1197), .B1(new_n1194), .B2(new_n1193), .C1(new_n1203), .C2(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1208), .A2(new_n723), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n778), .B1(G50), .B2(new_n1132), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n1179), .C2(new_n719), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1107), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1185), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n1126), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT115), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1110), .B2(new_n1123), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1102), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1179), .A2(new_n917), .A3(G330), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1170), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n917), .B2(G330), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n899), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1171), .A2(new_n1183), .A3(new_n1180), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1219), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n670), .B1(new_n1218), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1186), .B(new_n1212), .C1(new_n1214), .C2(new_n1227), .ZN(G375));
  INV_X1    g1028(.A(G303), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n990), .B1(new_n1229), .B2(new_n770), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n746), .A2(G294), .B1(new_n752), .B2(G107), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n455), .B2(new_n754), .C1(new_n814), .C2(new_n757), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n325), .B1(new_n979), .B2(new_n556), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1035), .A4(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n761), .A2(G50), .B1(G150), .B2(new_n752), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT122), .Z(new_n1236));
  OAI21_X1  g1036(.A(new_n1187), .B1(new_n1198), .B2(new_n770), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n749), .A2(G159), .B1(G137), .B2(new_n758), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n325), .B1(new_n755), .B2(new_n1134), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n800), .C2(new_n745), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n723), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n778), .C1(G68), .C2(new_n1132), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1087), .B2(new_n718), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1106), .B2(new_n960), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1103), .A2(new_n1109), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1247), .B2(new_n970), .ZN(G381));
  NAND2_X1  g1048(.A1(new_n1186), .A2(new_n1212), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n671), .B1(new_n1213), .B2(new_n1225), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1219), .B1(new_n1218), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G378), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G390), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1014), .A2(new_n782), .A3(new_n1047), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  OR4_X1    g1060(.A1(G387), .A2(new_n1255), .A3(G381), .A4(new_n1260), .ZN(G407));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G343), .C2(new_n1255), .ZN(G409));
  AND2_X1   g1062(.A1(new_n649), .A2(G213), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1211), .B1(new_n1264), .B2(new_n960), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1130), .A2(new_n1155), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1213), .A2(new_n969), .A3(new_n1185), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1263), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n671), .B1(new_n1246), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1247), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1245), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1257), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(G384), .A3(new_n1245), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1263), .A2(KEYINPUT123), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1263), .A2(G2897), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1268), .B(new_n1282), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT62), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G375), .A2(G378), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1268), .A4(new_n1282), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1281), .A2(new_n1284), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n782), .B1(new_n1014), .B2(new_n1047), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1259), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G390), .A2(new_n1005), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1004), .A2(new_n972), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n958), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n949), .A2(new_n953), .A3(new_n956), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n971), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1293), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1083), .A3(new_n1080), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G390), .A2(new_n1005), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1292), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT105), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1298), .A2(new_n1305), .ZN(new_n1306));
  AOI211_X1 g1106(.A(G390), .B(new_n1290), .C1(new_n1306), .C2(new_n1006), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT125), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(G390), .A2(new_n1290), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1302), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1310), .B(new_n1311), .C1(new_n1312), .C2(new_n1292), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1288), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1283), .A2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1268), .A4(new_n1282), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1281), .A2(new_n1317), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1315), .A2(KEYINPUT126), .A3(new_n1320), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(G405));
  NAND2_X1  g1125(.A1(new_n1285), .A2(new_n1255), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1282), .B(KEYINPUT127), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1326), .B(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1314), .ZN(G402));
endmodule


