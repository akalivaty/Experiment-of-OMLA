//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(G146), .C1(KEYINPUT16), .C2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT70), .B(G119), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n196), .A2(G128), .B1(KEYINPUT23), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n196), .B2(G128), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n202));
  INV_X1    g016(.A(G110), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(KEYINPUT70), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n197), .B2(G128), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT24), .B(G110), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(new_n201), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT79), .B1(new_n213), .B2(G110), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n195), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n193), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n192), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(G110), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n209), .A2(new_n210), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n187), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n205), .A2(new_n207), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT23), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n198), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n208), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n202), .B1(new_n229), .B2(new_n203), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n204), .A2(new_n211), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n194), .B(new_n192), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(KEYINPUT80), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G953), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(G221), .A3(G234), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT81), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G137), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n223), .A2(new_n234), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  OR3_X1    g057(.A1(new_n215), .A2(new_n222), .A3(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n242), .A2(KEYINPUT25), .A3(new_n243), .A4(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n243), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n242), .A2(new_n244), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(G902), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G472), .A2(G902), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(KEYINPUT32), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n260));
  NOR2_X1   g074(.A1(G237), .A2(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G210), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n260), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n193), .A2(G143), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT66), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT0), .A4(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT11), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(G137), .ZN(new_n279));
  INV_X1    g093(.A(G137), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT11), .A3(G134), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(G137), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  AOI21_X1  g098(.A(G131), .B1(new_n278), .B2(G137), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n268), .A2(G146), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n193), .A2(G143), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n271), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT0), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n225), .A3(KEYINPUT64), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT64), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(KEYINPUT0), .B2(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n290), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n293), .A2(new_n295), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n267), .A2(new_n269), .B1(KEYINPUT0), .B2(G128), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT65), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n276), .B(new_n287), .C1(new_n297), .C2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n205), .A2(new_n207), .A3(G116), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n303));
  INV_X1    g117(.A(G116), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT71), .A2(G116), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(G119), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT2), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G113), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n302), .A2(new_n307), .A3(new_n313), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n320));
  OAI22_X1  g134(.A1(new_n320), .A2(new_n269), .B1(new_n267), .B2(G128), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT68), .B1(new_n273), .B2(new_n320), .ZN(new_n323));
  AND4_X1   g137(.A1(KEYINPUT68), .A2(new_n320), .A3(new_n267), .A4(new_n269), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n279), .A2(new_n285), .A3(new_n281), .ZN(new_n326));
  INV_X1    g140(.A(G131), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n280), .A2(G134), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(new_n282), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n301), .A2(new_n319), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n266), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n301), .A2(KEYINPUT30), .A3(new_n331), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n301), .A2(new_n331), .A3(KEYINPUT72), .A4(KEYINPUT30), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n329), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT67), .A3(new_n286), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n326), .B2(new_n329), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n325), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n301), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n319), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n333), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT31), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT74), .B1(new_n347), .B2(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n317), .A2(new_n318), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(KEYINPUT75), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n332), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n319), .B1(new_n301), .B2(new_n343), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT28), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n332), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n266), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n349), .A2(new_n350), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n347), .A2(new_n348), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n291), .B1(new_n290), .B2(new_n296), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT65), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n364), .A2(new_n365), .B1(new_n272), .B2(new_n275), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n366), .A2(new_n287), .B1(new_n325), .B2(new_n330), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n354), .A2(KEYINPUT75), .B1(new_n367), .B2(new_n319), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n344), .A2(new_n351), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n357), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n358), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n360), .B(new_n265), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n259), .B1(new_n361), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n356), .A2(new_n377), .A3(new_n358), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n301), .A2(new_n331), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n351), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n357), .B1(new_n381), .B2(new_n332), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n379), .B(KEYINPUT29), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n266), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n332), .ZN(new_n386));
  AOI211_X1 g200(.A(new_n386), .B(new_n266), .C1(new_n338), .C2(new_n346), .ZN(new_n387));
  AOI21_X1  g201(.A(G902), .B1(new_n387), .B2(new_n377), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G472), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT77), .B(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n338), .A2(new_n346), .ZN(new_n393));
  INV_X1    g207(.A(new_n333), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n348), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n348), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n265), .B1(new_n372), .B2(new_n373), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT76), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n399), .A2(new_n401), .A3(new_n363), .A4(new_n374), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n392), .B1(new_n402), .B2(new_n258), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n257), .B1(new_n391), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n258), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n397), .A2(new_n398), .B1(new_n400), .B2(KEYINPUT76), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n362), .B1(new_n359), .B2(new_n360), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n376), .B(new_n390), .C1(new_n410), .C2(new_n392), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT83), .A3(new_n257), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT84), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n250), .A2(G953), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n225), .A2(G143), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n225), .A2(G143), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(KEYINPUT13), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n278), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n268), .A2(G128), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT13), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT91), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(new_n423), .A3(new_n278), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n427), .B(KEYINPUT92), .Z(new_n428));
  NAND3_X1  g242(.A1(new_n305), .A2(G122), .A3(new_n306), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n304), .A2(G122), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G107), .ZN(new_n432));
  INV_X1    g246(.A(G107), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n426), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n419), .ZN(new_n437));
  OAI21_X1  g251(.A(G134), .B1(new_n437), .B2(new_n418), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n427), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n434), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT14), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(new_n429), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT93), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n433), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n429), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT93), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n440), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n416), .B(new_n417), .C1(new_n436), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n448), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n439), .A2(new_n434), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n416), .A2(new_n417), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n426), .A2(new_n428), .A3(new_n435), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n243), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n450), .A2(new_n243), .A3(new_n456), .A4(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(KEYINPUT94), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT94), .B1(new_n460), .B2(new_n462), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G104), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(G104), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT90), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n261), .A2(G143), .A3(G214), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G143), .B1(new_n261), .B2(G214), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT18), .B(G131), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G125), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G140), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n191), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G146), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n194), .ZN(new_n481));
  INV_X1    g295(.A(new_n475), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n327), .A3(new_n473), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n218), .B(new_n192), .C1(new_n488), .C2(new_n486), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n472), .B(new_n485), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n490), .A2(new_n489), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n471), .B1(new_n493), .B2(new_n485), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n243), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G475), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n235), .A2(G952), .ZN(new_n497));
  INV_X1    g311(.A(G234), .ZN(new_n498));
  INV_X1    g312(.A(G237), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n243), .B(new_n235), .C1(G234), .C2(G237), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT21), .B(G898), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n479), .B(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n192), .B1(new_n507), .B2(G146), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n486), .A2(new_n487), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n485), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n470), .B2(new_n469), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n491), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(G475), .A2(G902), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n506), .A3(new_n513), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n496), .B(new_n505), .C1(new_n514), .C2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n414), .B1(new_n466), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n465), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n463), .ZN(new_n520));
  INV_X1    g334(.A(new_n514), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n521), .A2(new_n515), .B1(G475), .B2(new_n495), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n520), .A2(KEYINPUT95), .A3(new_n505), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G214), .B1(G237), .B2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G210), .B1(G237), .B2(G902), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT6), .ZN(new_n530));
  INV_X1    g344(.A(G104), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT3), .B1(new_n531), .B2(G107), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT3), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n433), .A3(G104), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(G107), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT4), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n536), .A2(new_n537), .A3(G101), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n317), .B2(new_n318), .ZN(new_n539));
  AOI21_X1  g353(.A(G101), .B1(new_n531), .B2(G107), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n540), .A3(new_n534), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT85), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n532), .A2(new_n540), .A3(new_n534), .A4(KEYINPUT85), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n537), .B1(new_n536), .B2(G101), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n302), .A2(new_n307), .A3(KEYINPUT5), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT5), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n205), .A2(new_n207), .A3(new_n549), .A4(G116), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n550), .A2(G113), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n302), .A2(new_n307), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n548), .A2(new_n551), .B1(new_n552), .B2(new_n313), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n433), .A2(G104), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n535), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n555), .A2(G101), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n543), .B2(new_n544), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n539), .A2(new_n547), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G122), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n530), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n558), .B2(KEYINPUT88), .ZN(new_n562));
  INV_X1    g376(.A(new_n538), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n547), .A2(new_n351), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n557), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT88), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n529), .B(new_n560), .C1(new_n562), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n565), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n530), .A4(new_n561), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n561), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n529), .B1(new_n574), .B2(new_n560), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n366), .A2(new_n477), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n325), .A2(G125), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G224), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G953), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n578), .B(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n573), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n578), .ZN(new_n583));
  INV_X1    g397(.A(new_n580), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT7), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n553), .B(new_n557), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n559), .B(KEYINPUT8), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n583), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n585), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n578), .A2(new_n589), .B1(new_n558), .B2(new_n559), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n528), .B1(new_n582), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n560), .B1(new_n562), .B2(new_n566), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT89), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n578), .B(new_n584), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n572), .A3(new_n567), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n591), .A3(new_n527), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n526), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n416), .A2(new_n243), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n600), .A2(G221), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n321), .A2(KEYINPUT86), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT86), .ZN(new_n603));
  OAI221_X1 g417(.A(new_n603), .B1(new_n267), .B2(G128), .C1(new_n269), .C2(new_n320), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n602), .B(new_n604), .C1(new_n323), .C2(new_n324), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n557), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n366), .A2(new_n547), .A3(new_n563), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n557), .A2(new_n325), .A3(KEYINPUT10), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT87), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT87), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n608), .A2(new_n609), .A3(new_n613), .A4(new_n610), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n287), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n287), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n608), .A2(new_n609), .A3(new_n616), .A4(new_n610), .ZN(new_n617));
  XNOR2_X1  g431(.A(G110), .B(G140), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n235), .A2(G227), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n618), .B(new_n619), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n556), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n545), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n273), .A2(new_n320), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT68), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n320), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n321), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n606), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT12), .B1(new_n632), .B2(new_n287), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT12), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n634), .B(new_n616), .C1(new_n631), .C2(new_n606), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n617), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n615), .A2(new_n623), .B1(new_n636), .B2(new_n620), .ZN(new_n637));
  OAI21_X1  g451(.A(G469), .B1(new_n637), .B2(G902), .ZN(new_n638));
  INV_X1    g452(.A(G469), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n621), .B1(new_n615), .B2(new_n617), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n633), .A2(new_n635), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n622), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n639), .B(new_n243), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n601), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n524), .A2(new_n599), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n413), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G101), .ZN(G3));
  OAI21_X1  g462(.A(new_n243), .B1(new_n361), .B2(new_n375), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n649), .A2(G472), .B1(new_n258), .B2(new_n402), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n638), .A2(new_n643), .ZN(new_n651));
  INV_X1    g465(.A(new_n601), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n256), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n597), .A2(new_n591), .A3(new_n527), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n527), .B1(new_n597), .B2(new_n591), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n505), .B(new_n525), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n457), .A2(new_n458), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n660), .B(new_n454), .C1(new_n436), .C2(new_n449), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n454), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n453), .A2(new_n455), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(KEYINPUT33), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT97), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(KEYINPUT97), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n450), .A2(new_n456), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n665), .B(new_n666), .C1(KEYINPUT33), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n243), .A2(G478), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n659), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n496), .B1(new_n516), .B2(new_n514), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n658), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n655), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n531), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n466), .A2(new_n522), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n658), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n679), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n599), .A2(KEYINPUT99), .A3(new_n505), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n655), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT35), .B(G107), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  OAI21_X1  g500(.A(new_n525), .B1(new_n656), .B2(new_n657), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n653), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n524), .A3(new_n650), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n223), .A2(new_n234), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n223), .B(new_n234), .C1(KEYINPUT36), .C2(new_n241), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n693), .A2(new_n254), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT100), .B1(new_n252), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n251), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n247), .B2(new_n248), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n695), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n690), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n252), .A2(KEYINPUT100), .A3(new_n696), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n700), .B1(new_n699), .B2(new_n695), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(KEYINPUT101), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n689), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT37), .B(G110), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT102), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n707), .B(new_n709), .ZN(G12));
  AND3_X1   g524(.A1(new_n703), .A2(KEYINPUT101), .A3(new_n704), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT101), .B1(new_n703), .B2(new_n704), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n644), .B(new_n525), .C1(new_n657), .C2(new_n656), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n258), .B1(new_n361), .B2(new_n375), .ZN(new_n715));
  INV_X1    g529(.A(new_n392), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n402), .A2(new_n259), .B1(G472), .B2(new_n389), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(G900), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n502), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n500), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n679), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n713), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G128), .ZN(G30));
  NAND2_X1  g540(.A1(new_n593), .A2(new_n598), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n703), .A2(new_n704), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n525), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n466), .A2(new_n671), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n393), .A2(new_n332), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n266), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n381), .A2(new_n332), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n737), .B(new_n243), .C1(new_n266), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G472), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n376), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n735), .B1(new_n741), .B2(new_n403), .ZN(new_n742));
  OR3_X1    g556(.A1(new_n732), .A2(new_n733), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n733), .B1(new_n732), .B2(new_n742), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n722), .B(KEYINPUT39), .Z(new_n745));
  OR2_X1    g559(.A1(new_n653), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT40), .Z(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT105), .B(G143), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G45));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n670), .A2(new_n671), .A3(new_n722), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n713), .A2(new_n719), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n688), .A2(new_n411), .A3(new_n752), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT106), .B1(new_n754), .B2(new_n706), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G146), .ZN(G48));
  OAI21_X1  g571(.A(new_n243), .B1(new_n640), .B2(new_n642), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(G469), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n652), .A3(new_n643), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n404), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n673), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT41), .B(G113), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n683), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G116), .ZN(G18));
  INV_X1    g580(.A(new_n760), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n524), .A2(new_n599), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n713), .A2(new_n411), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT107), .B(G119), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G21));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n379), .B(new_n265), .C1(new_n382), .C2(new_n383), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n363), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n773), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT108), .B1(new_n775), .B2(new_n362), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n776), .A3(new_n399), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n649), .A2(G472), .B1(new_n777), .B2(new_n258), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(new_n257), .ZN(new_n779));
  INV_X1    g593(.A(new_n658), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n760), .A2(new_n734), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G122), .ZN(G24));
  NOR2_X1   g597(.A1(new_n687), .A2(new_n760), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n778), .A3(new_n730), .A4(new_n752), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G125), .ZN(G27));
  AOI21_X1  g600(.A(KEYINPUT32), .B1(new_n402), .B2(new_n258), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n752), .B(new_n257), .C1(new_n391), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n653), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n644), .A2(KEYINPUT109), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n656), .A2(new_n657), .A3(new_n526), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT42), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n644), .A2(KEYINPUT109), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n789), .B(new_n601), .C1(new_n638), .C2(new_n643), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n593), .A2(new_n525), .A3(new_n598), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n256), .B1(new_n717), .B2(new_n718), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n752), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n327), .ZN(G33));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n799), .A3(new_n724), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NAND2_X1  g619(.A1(new_n670), .A2(new_n522), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT43), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n650), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n730), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n637), .A2(KEYINPUT45), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n637), .A2(KEYINPUT45), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(G469), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(G469), .A2(G902), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT46), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n815), .A2(KEYINPUT46), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n643), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n652), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n745), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n811), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n812), .A2(new_n792), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G137), .ZN(G39));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n822), .B(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n752), .A2(new_n792), .A3(new_n256), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n411), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  NAND4_X1  g646(.A1(new_n762), .A2(new_n765), .A3(new_n769), .A4(new_n782), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n802), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n460), .A2(new_n462), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n671), .A2(new_n836), .A3(KEYINPUT111), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT111), .B1(new_n671), .B2(new_n836), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n672), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n780), .A2(new_n650), .A3(new_n839), .A4(new_n654), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n689), .B2(new_n706), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n647), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n798), .A2(new_n730), .A3(new_n752), .A4(new_n778), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n522), .A2(new_n836), .A3(new_n722), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n797), .A2(new_n653), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n702), .A3(new_n411), .A4(new_n705), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n844), .A2(new_n804), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n688), .A2(new_n411), .A3(new_n724), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n785), .B1(new_n850), .B2(new_n706), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n699), .A2(new_n695), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT112), .B1(new_n852), .B2(new_n722), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n699), .A2(new_n695), .A3(new_n854), .A4(new_n723), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n742), .A2(new_n856), .A3(new_n714), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n858), .A2(new_n756), .A3(KEYINPUT52), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n858), .B2(new_n756), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n834), .B(new_n849), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n753), .A2(new_n755), .ZN(new_n865));
  INV_X1    g679(.A(new_n742), .ZN(new_n866));
  INV_X1    g680(.A(new_n856), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n688), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n725), .A3(new_n785), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n864), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n858), .A2(new_n756), .A3(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n411), .A2(new_n257), .A3(new_n767), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n680), .B2(new_n682), .ZN(new_n874));
  INV_X1    g688(.A(new_n673), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n778), .A2(new_n257), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n781), .A2(new_n505), .A3(new_n599), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n873), .A2(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n794), .A2(new_n801), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n769), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n645), .B1(new_n406), .B2(new_n412), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n841), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n844), .A2(new_n804), .A3(new_n847), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n872), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT54), .B1(new_n863), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n861), .A2(new_n862), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n848), .A2(new_n882), .A3(new_n841), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT113), .B1(new_n883), .B2(new_n884), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n833), .A2(new_n862), .A3(new_n802), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n872), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n889), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n779), .A2(new_n501), .A3(new_n808), .ZN(new_n899));
  INV_X1    g713(.A(new_n729), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n526), .A3(new_n767), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(KEYINPUT50), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n902), .B(new_n904), .Z(new_n905));
  OR3_X1    g719(.A1(new_n899), .A2(KEYINPUT114), .A3(new_n797), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT114), .B1(new_n899), .B2(new_n797), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n759), .A2(new_n643), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(new_n652), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n906), .B(new_n907), .C1(new_n828), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n741), .A2(new_n403), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n797), .A2(new_n760), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(new_n501), .A3(new_n257), .A4(new_n912), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n671), .A3(new_n670), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n807), .A2(new_n500), .A3(new_n760), .A4(new_n797), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n778), .A2(new_n730), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n905), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n905), .A2(KEYINPUT51), .A3(new_n910), .A4(new_n917), .ZN(new_n921));
  INV_X1    g735(.A(new_n787), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n256), .B1(new_n922), .B2(new_n718), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT48), .Z(new_n925));
  INV_X1    g739(.A(new_n784), .ZN(new_n926));
  OAI221_X1 g740(.A(new_n497), .B1(new_n672), .B2(new_n913), .C1(new_n899), .C2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n920), .A2(new_n921), .A3(new_n928), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n898), .A2(new_n929), .B1(G952), .B2(G953), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n256), .A2(new_n526), .A3(new_n601), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT110), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n522), .B(new_n670), .C1(new_n908), .C2(KEYINPUT49), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(KEYINPUT49), .B2(new_n908), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n932), .A2(new_n911), .A3(new_n900), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT116), .ZN(G75));
  NAND4_X1  g751(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT53), .A4(new_n769), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n870), .B2(new_n871), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n862), .A2(new_n861), .B1(new_n939), .B2(new_n893), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n243), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(G210), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n595), .A2(new_n572), .A3(new_n567), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n596), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n942), .B2(new_n943), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n235), .A2(G952), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G51));
  NOR3_X1   g764(.A1(new_n940), .A2(new_n243), .A3(new_n815), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n816), .B(KEYINPUT57), .Z(new_n952));
  OAI21_X1  g766(.A(new_n894), .B1(new_n859), .B2(new_n860), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n885), .A2(new_n890), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT113), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT54), .B1(new_n957), .B2(new_n887), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n889), .A2(new_n895), .A3(KEYINPUT117), .A4(new_n896), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT117), .B1(new_n940), .B2(new_n896), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n640), .A2(new_n642), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT118), .Z(new_n964));
  AOI21_X1  g778(.A(new_n951), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT119), .B1(new_n965), .B2(new_n949), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT119), .ZN(new_n967));
  INV_X1    g781(.A(new_n949), .ZN(new_n968));
  INV_X1    g782(.A(new_n964), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT117), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n897), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n958), .A3(new_n959), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n972), .B2(new_n952), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n967), .B(new_n968), .C1(new_n973), .C2(new_n951), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n966), .A2(new_n974), .ZN(G54));
  NAND3_X1  g789(.A1(new_n941), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  INV_X1    g790(.A(new_n512), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n976), .A2(KEYINPUT120), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT120), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(G60));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT59), .Z(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n888), .B2(new_n897), .ZN(new_n984));
  INV_X1    g798(.A(new_n668), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n968), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n668), .A2(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n972), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT121), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT121), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(G63));
  NAND2_X1  g805(.A1(G217), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT60), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n940), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n693), .A3(new_n694), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n995), .B(new_n968), .C1(new_n253), .C2(new_n994), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G66));
  OAI21_X1  g812(.A(G953), .B1(new_n503), .B2(new_n579), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT122), .Z(new_n1000));
  NOR2_X1   g814(.A1(new_n843), .A2(new_n833), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT123), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n944), .B1(G898), .B2(new_n235), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  NAND2_X1  g819(.A1(new_n344), .A2(new_n345), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n338), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT124), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(new_n507), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G900), .A2(G953), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n823), .A2(new_n599), .A3(new_n735), .A4(new_n923), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1011), .A2(new_n880), .A3(new_n804), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n865), .A2(new_n851), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n825), .A3(new_n831), .A4(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1009), .B(new_n1010), .C1(new_n1014), .C2(G953), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n235), .B1(G227), .B2(G900), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT126), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT62), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1013), .A2(new_n748), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT125), .Z(new_n1020));
  INV_X1    g834(.A(new_n746), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n413), .A2(new_n1021), .A3(new_n792), .A4(new_n839), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n825), .A2(new_n831), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1018), .B1(new_n1013), .B2(new_n748), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(G953), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1015), .B(new_n1017), .C1(new_n1026), .C2(new_n1009), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1027), .A2(KEYINPUT127), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1027), .A2(KEYINPUT127), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1015), .B1(new_n1026), .B2(new_n1009), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n1016), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1028), .B1(new_n1029), .B2(new_n1031), .ZN(G72));
  NAND3_X1  g846(.A1(new_n1020), .A2(new_n1001), .A3(new_n1025), .ZN(new_n1033));
  NAND2_X1  g847(.A1(G472), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT63), .Z(new_n1035));
  AOI21_X1  g849(.A(new_n737), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n863), .A2(new_n887), .ZN(new_n1037));
  INV_X1    g851(.A(new_n387), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1038), .A2(new_n737), .A3(new_n1035), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1001), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1035), .B1(new_n1014), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n1042), .A2(new_n387), .ZN(new_n1043));
  NOR4_X1   g857(.A1(new_n1036), .A2(new_n949), .A3(new_n1040), .A4(new_n1043), .ZN(G57));
endmodule


