

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(n704), .B(KEYINPUT90), .ZN(n773) );
  NAND2_X1 U555 ( .A1(n703), .A2(n807), .ZN(n747) );
  NOR2_X1 U556 ( .A1(n521), .A2(n531), .ZN(n529) );
  INV_X1 U557 ( .A(n532), .ZN(n531) );
  XNOR2_X1 U558 ( .A(n747), .B(KEYINPUT93), .ZN(n732) );
  NAND2_X1 U559 ( .A1(n731), .A2(n544), .ZN(n543) );
  INV_X1 U560 ( .A(n980), .ZN(n544) );
  NOR2_X1 U561 ( .A1(n819), .A2(n523), .ZN(n532) );
  XNOR2_X1 U562 ( .A(n542), .B(KEYINPUT96), .ZN(n736) );
  NAND2_X1 U563 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U564 ( .A1(n543), .A2(n986), .ZN(n540) );
  NAND2_X1 U565 ( .A1(n525), .A2(n746), .ZN(n760) );
  XNOR2_X1 U566 ( .A(n745), .B(n526), .ZN(n525) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n526) );
  INV_X1 U568 ( .A(KEYINPUT98), .ZN(n539) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n807) );
  NAND2_X1 U570 ( .A1(n552), .A2(n534), .ZN(n533) );
  INV_X1 U571 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U572 ( .A1(n787), .A2(n532), .ZN(n530) );
  NOR2_X1 U573 ( .A1(n529), .A2(n520), .ZN(n528) );
  NOR2_X1 U574 ( .A1(n556), .A2(n555), .ZN(G160) );
  XNOR2_X1 U575 ( .A(KEYINPUT101), .B(n831), .ZN(n520) );
  AND2_X1 U576 ( .A1(n786), .A2(n545), .ZN(n521) );
  XOR2_X1 U577 ( .A(KEYINPUT84), .B(n559), .Z(n522) );
  AND2_X1 U578 ( .A1(n988), .A2(n830), .ZN(n523) );
  XOR2_X1 U579 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n524) );
  NAND2_X1 U580 ( .A1(n527), .A2(n760), .ZN(n757) );
  AND2_X1 U581 ( .A1(n759), .A2(n753), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n530), .A2(n528), .ZN(n832) );
  NAND2_X1 U583 ( .A1(n905), .A2(G138), .ZN(n558) );
  XNOR2_X2 U584 ( .A(n533), .B(KEYINPUT17), .ZN(n905) );
  INV_X1 U585 ( .A(n538), .ZN(n783) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U587 ( .A(n767), .B(n539), .ZN(n535) );
  XNOR2_X1 U588 ( .A(n758), .B(n524), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n990), .ZN(n769) );
  NAND2_X1 U590 ( .A1(n538), .A2(n991), .ZN(n537) );
  OR2_X1 U591 ( .A1(n730), .A2(n543), .ZN(n737) );
  INV_X1 U592 ( .A(n730), .ZN(n541) );
  OR2_X1 U593 ( .A1(n785), .A2(n784), .ZN(n545) );
  INV_X1 U594 ( .A(KEYINPUT30), .ZN(n708) );
  XNOR2_X1 U595 ( .A(n708), .B(KEYINPUT97), .ZN(n709) );
  XNOR2_X1 U596 ( .A(n710), .B(n709), .ZN(n711) );
  INV_X1 U597 ( .A(KEYINPUT31), .ZN(n719) );
  INV_X1 U598 ( .A(n982), .ZN(n776) );
  NAND2_X1 U599 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U600 ( .A1(n644), .A2(G651), .ZN(n673) );
  AND2_X1 U601 ( .A1(G2104), .A2(G2105), .ZN(n901) );
  NAND2_X1 U602 ( .A1(G113), .A2(n901), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT66), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G137), .A2(n905), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT67), .B(n547), .Z(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n556) );
  INV_X1 U607 ( .A(G2104), .ZN(n552) );
  NOR2_X2 U608 ( .A1(G2105), .A2(n552), .ZN(n622) );
  NAND2_X1 U609 ( .A1(G101), .A2(n622), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT65), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT23), .ZN(n554) );
  AND2_X1 U612 ( .A1(n552), .A2(G2105), .ZN(n900) );
  NAND2_X1 U613 ( .A1(G125), .A2(n900), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G102), .A2(n622), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n901), .A2(G114), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n522), .A2(n560), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G126), .A2(n900), .ZN(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT83), .B(n561), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G164) );
  INV_X1 U622 ( .A(G651), .ZN(n567) );
  NOR2_X1 U623 ( .A1(G543), .A2(n567), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT1), .B(n564), .Z(n664) );
  NAND2_X1 U625 ( .A1(G64), .A2(n664), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  NAND2_X1 U627 ( .A1(G52), .A2(n673), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n572) );
  NOR2_X1 U629 ( .A1(G543), .A2(G651), .ZN(n665) );
  NAND2_X1 U630 ( .A1(G90), .A2(n665), .ZN(n569) );
  NOR2_X1 U631 ( .A1(n644), .A2(n567), .ZN(n668) );
  NAND2_X1 U632 ( .A1(G77), .A2(n668), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U635 ( .A1(n572), .A2(n571), .ZN(G171) );
  AND2_X1 U636 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U637 ( .A(G132), .ZN(G219) );
  INV_X1 U638 ( .A(G82), .ZN(G220) );
  INV_X1 U639 ( .A(G57), .ZN(G237) );
  NAND2_X1 U640 ( .A1(n665), .A2(G89), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G76), .A2(n668), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT5), .B(n576), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G63), .A2(n664), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G51), .A2(n673), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT6), .B(KEYINPUT72), .Z(n579) );
  XNOR2_X1 U649 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U651 ( .A(KEYINPUT7), .B(n583), .ZN(G168) );
  XOR2_X1 U652 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n833) );
  NAND2_X1 U656 ( .A1(n833), .A2(G567), .ZN(n585) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U658 ( .A1(G56), .A2(n664), .ZN(n586) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n586), .Z(n592) );
  NAND2_X1 U660 ( .A1(n665), .A2(G81), .ZN(n587) );
  XNOR2_X1 U661 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G68), .A2(n668), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n673), .A2(G43), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n980) );
  INV_X1 U668 ( .A(G860), .ZN(n633) );
  NOR2_X1 U669 ( .A1(n980), .A2(n633), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT70), .B(n595), .Z(G153) );
  INV_X1 U671 ( .A(G868), .ZN(n684) );
  NOR2_X1 U672 ( .A1(n684), .A2(G171), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n596), .B(KEYINPUT71), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G79), .A2(n668), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G54), .A2(n673), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U677 ( .A1(G66), .A2(n664), .ZN(n600) );
  NAND2_X1 U678 ( .A1(G92), .A2(n665), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT15), .ZN(n986) );
  NAND2_X1 U682 ( .A1(n684), .A2(n986), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U684 ( .A1(G65), .A2(n664), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G53), .A2(n673), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U687 ( .A(KEYINPUT69), .B(n608), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G91), .A2(n665), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G78), .A2(n668), .ZN(n609) );
  AND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(G299) );
  INV_X1 U692 ( .A(G299), .ZN(n996) );
  NAND2_X1 U693 ( .A1(n996), .A2(n684), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n613), .B(KEYINPUT73), .ZN(n615) );
  NOR2_X1 U695 ( .A1(n684), .A2(G286), .ZN(n614) );
  NOR2_X1 U696 ( .A1(n615), .A2(n614), .ZN(G297) );
  NAND2_X1 U697 ( .A1(n633), .A2(G559), .ZN(n616) );
  INV_X1 U698 ( .A(n986), .ZN(n631) );
  NAND2_X1 U699 ( .A1(n616), .A2(n631), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U701 ( .A1(G868), .A2(n980), .ZN(n620) );
  NAND2_X1 U702 ( .A1(G868), .A2(n631), .ZN(n618) );
  NOR2_X1 U703 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U704 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U705 ( .A1(n900), .A2(G123), .ZN(n621) );
  XNOR2_X1 U706 ( .A(n621), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G99), .A2(n622), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G111), .A2(n901), .ZN(n626) );
  NAND2_X1 U710 ( .A1(G135), .A2(n905), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n930) );
  XNOR2_X1 U713 ( .A(n930), .B(G2096), .ZN(n630) );
  INV_X1 U714 ( .A(G2100), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U716 ( .A1(G559), .A2(n631), .ZN(n632) );
  XOR2_X1 U717 ( .A(n980), .B(n632), .Z(n682) );
  NAND2_X1 U718 ( .A1(n633), .A2(n682), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G80), .A2(n668), .ZN(n634) );
  XNOR2_X1 U720 ( .A(n634), .B(KEYINPUT74), .ZN(n641) );
  NAND2_X1 U721 ( .A1(G67), .A2(n664), .ZN(n636) );
  NAND2_X1 U722 ( .A1(G93), .A2(n665), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G55), .A2(n673), .ZN(n637) );
  XNOR2_X1 U725 ( .A(KEYINPUT75), .B(n637), .ZN(n638) );
  NOR2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n685) );
  XNOR2_X1 U728 ( .A(n642), .B(n685), .ZN(G145) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n643) );
  XNOR2_X1 U730 ( .A(n643), .B(KEYINPUT76), .ZN(n649) );
  NAND2_X1 U731 ( .A1(G49), .A2(n673), .ZN(n646) );
  NAND2_X1 U732 ( .A1(G87), .A2(n644), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U734 ( .A1(n664), .A2(n647), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U736 ( .A1(G85), .A2(n665), .ZN(n651) );
  NAND2_X1 U737 ( .A1(G72), .A2(n668), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U739 ( .A1(G60), .A2(n664), .ZN(n653) );
  NAND2_X1 U740 ( .A1(G47), .A2(n673), .ZN(n652) );
  NAND2_X1 U741 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U742 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U743 ( .A(KEYINPUT68), .B(n656), .Z(G290) );
  NAND2_X1 U744 ( .A1(G62), .A2(n664), .ZN(n658) );
  NAND2_X1 U745 ( .A1(G88), .A2(n665), .ZN(n657) );
  NAND2_X1 U746 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n668), .A2(G75), .ZN(n659) );
  XOR2_X1 U748 ( .A(KEYINPUT78), .B(n659), .Z(n660) );
  NOR2_X1 U749 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n673), .A2(G50), .ZN(n662) );
  NAND2_X1 U751 ( .A1(n663), .A2(n662), .ZN(G303) );
  INV_X1 U752 ( .A(G303), .ZN(G166) );
  NAND2_X1 U753 ( .A1(G61), .A2(n664), .ZN(n667) );
  NAND2_X1 U754 ( .A1(G86), .A2(n665), .ZN(n666) );
  NAND2_X1 U755 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U756 ( .A1(n668), .A2(G73), .ZN(n669) );
  XOR2_X1 U757 ( .A(KEYINPUT2), .B(n669), .Z(n670) );
  NOR2_X1 U758 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U759 ( .A(KEYINPUT77), .B(n672), .Z(n675) );
  NAND2_X1 U760 ( .A1(n673), .A2(G48), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(G305) );
  XOR2_X1 U762 ( .A(KEYINPUT19), .B(KEYINPUT79), .Z(n676) );
  XNOR2_X1 U763 ( .A(G288), .B(n676), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n685), .B(n677), .ZN(n679) );
  XNOR2_X1 U765 ( .A(G290), .B(G166), .ZN(n678) );
  XNOR2_X1 U766 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n680), .B(G305), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n681), .B(G299), .ZN(n915) );
  XOR2_X1 U769 ( .A(n915), .B(n682), .Z(n683) );
  NOR2_X1 U770 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U771 ( .A1(G868), .A2(n685), .ZN(n686) );
  NOR2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U773 ( .A(KEYINPUT80), .B(n688), .ZN(G295) );
  NAND2_X1 U774 ( .A1(G2078), .A2(G2084), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT20), .B(n689), .Z(n690) );
  NAND2_X1 U776 ( .A1(G2090), .A2(n690), .ZN(n691) );
  XNOR2_X1 U777 ( .A(KEYINPUT21), .B(n691), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n692), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U779 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U780 ( .A1(G69), .A2(G120), .ZN(n693) );
  NOR2_X1 U781 ( .A1(G237), .A2(n693), .ZN(n694) );
  NAND2_X1 U782 ( .A1(G108), .A2(n694), .ZN(n927) );
  NAND2_X1 U783 ( .A1(n927), .A2(G567), .ZN(n701) );
  NOR2_X1 U784 ( .A1(G220), .A2(G219), .ZN(n695) );
  XOR2_X1 U785 ( .A(KEYINPUT22), .B(n695), .Z(n696) );
  NOR2_X1 U786 ( .A1(G218), .A2(n696), .ZN(n697) );
  XOR2_X1 U787 ( .A(KEYINPUT81), .B(n697), .Z(n698) );
  NAND2_X1 U788 ( .A1(G96), .A2(n698), .ZN(n699) );
  XNOR2_X1 U789 ( .A(KEYINPUT82), .B(n699), .ZN(n926) );
  NAND2_X1 U790 ( .A1(G2106), .A2(n926), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n838) );
  NAND2_X1 U792 ( .A1(G661), .A2(G483), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n838), .A2(n702), .ZN(n837) );
  NAND2_X1 U794 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U795 ( .A1(G160), .A2(G40), .ZN(n806) );
  INV_X1 U796 ( .A(n806), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n747), .A2(G8), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n773), .A2(G1966), .ZN(n706) );
  INV_X1 U799 ( .A(KEYINPUT91), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n706), .B(n705), .ZN(n761) );
  NOR2_X1 U801 ( .A1(G2084), .A2(n747), .ZN(n762) );
  NOR2_X1 U802 ( .A1(n761), .A2(n762), .ZN(n707) );
  NAND2_X1 U803 ( .A1(G8), .A2(n707), .ZN(n710) );
  NOR2_X1 U804 ( .A1(G168), .A2(n711), .ZN(n718) );
  INV_X1 U805 ( .A(n747), .ZN(n727) );
  NOR2_X1 U806 ( .A1(n727), .A2(G1961), .ZN(n712) );
  XNOR2_X1 U807 ( .A(n712), .B(KEYINPUT92), .ZN(n715) );
  XOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .Z(n713) );
  XNOR2_X1 U809 ( .A(KEYINPUT94), .B(n713), .ZN(n957) );
  INV_X1 U810 ( .A(n732), .ZN(n723) );
  NOR2_X1 U811 ( .A1(n957), .A2(n723), .ZN(n714) );
  NOR2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U813 ( .A(KEYINPUT95), .B(n716), .ZN(n721) );
  NOR2_X1 U814 ( .A1(G171), .A2(n721), .ZN(n717) );
  NOR2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U816 ( .A(n720), .B(n719), .ZN(n759) );
  NAND2_X1 U817 ( .A1(n721), .A2(G171), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n732), .A2(G2072), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n722), .B(KEYINPUT27), .ZN(n725) );
  AND2_X1 U820 ( .A1(G1956), .A2(n723), .ZN(n724) );
  NOR2_X1 U821 ( .A1(n725), .A2(n724), .ZN(n740) );
  NOR2_X1 U822 ( .A1(n996), .A2(n740), .ZN(n726) );
  XOR2_X1 U823 ( .A(n726), .B(KEYINPUT28), .Z(n744) );
  XOR2_X1 U824 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n729) );
  NAND2_X1 U825 ( .A1(n727), .A2(G1996), .ZN(n728) );
  XNOR2_X1 U826 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U827 ( .A1(G1341), .A2(n747), .ZN(n731) );
  NAND2_X1 U828 ( .A1(G1348), .A2(n747), .ZN(n734) );
  NAND2_X1 U829 ( .A1(G2067), .A2(n732), .ZN(n733) );
  NAND2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n737), .A2(n986), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n996), .A2(n740), .ZN(n741) );
  NAND2_X1 U835 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  INV_X1 U837 ( .A(G8), .ZN(n752) );
  NOR2_X1 U838 ( .A1(n773), .A2(G1971), .ZN(n749) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n750), .A2(G303), .ZN(n751) );
  OR2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  INV_X1 U843 ( .A(n753), .ZN(n755) );
  AND2_X1 U844 ( .A1(G286), .A2(G8), .ZN(n754) );
  OR2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n766) );
  INV_X1 U848 ( .A(n761), .ZN(n764) );
  NAND2_X1 U849 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n772) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n768) );
  NOR2_X1 U854 ( .A1(n772), .A2(n768), .ZN(n991) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n990) );
  XNOR2_X1 U856 ( .A(n769), .B(KEYINPUT100), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n770), .A2(n773), .ZN(n771) );
  NOR2_X1 U858 ( .A1(KEYINPUT33), .A2(n771), .ZN(n778) );
  XNOR2_X1 U859 ( .A(G1981), .B(G305), .ZN(n982) );
  AND2_X1 U860 ( .A1(n772), .A2(KEYINPUT33), .ZN(n774) );
  INV_X1 U861 ( .A(n773), .ZN(n784) );
  NAND2_X1 U862 ( .A1(n774), .A2(n784), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n787) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(KEYINPUT24), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n780), .A2(n784), .ZN(n786) );
  NAND2_X1 U867 ( .A1(G166), .A2(G8), .ZN(n781) );
  NOR2_X1 U868 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n785) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(KEYINPUT86), .Z(n789) );
  NAND2_X1 U871 ( .A1(G105), .A2(n622), .ZN(n788) );
  XNOR2_X1 U872 ( .A(n789), .B(n788), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G129), .A2(n900), .ZN(n791) );
  NAND2_X1 U874 ( .A1(G141), .A2(n905), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U877 ( .A1(n901), .A2(G117), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n795), .A2(n794), .ZN(n891) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n891), .ZN(n796) );
  XOR2_X1 U880 ( .A(KEYINPUT87), .B(n796), .Z(n805) );
  NAND2_X1 U881 ( .A1(G119), .A2(n900), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G95), .A2(n622), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G131), .A2(n905), .ZN(n799) );
  XNOR2_X1 U885 ( .A(KEYINPUT85), .B(n799), .ZN(n800) );
  NOR2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n901), .A2(G107), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n888) );
  NAND2_X1 U889 ( .A1(G1991), .A2(n888), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n805), .A2(n804), .ZN(n931) );
  NOR2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n830) );
  NAND2_X1 U892 ( .A1(n931), .A2(n830), .ZN(n808) );
  XOR2_X1 U893 ( .A(KEYINPUT88), .B(n808), .Z(n822) );
  XNOR2_X1 U894 ( .A(KEYINPUT89), .B(n822), .ZN(n818) );
  NAND2_X1 U895 ( .A1(G140), .A2(n905), .ZN(n810) );
  NAND2_X1 U896 ( .A1(G104), .A2(n622), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n811), .ZN(n816) );
  NAND2_X1 U899 ( .A1(G128), .A2(n900), .ZN(n813) );
  NAND2_X1 U900 ( .A1(G116), .A2(n901), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U903 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U904 ( .A(KEYINPUT36), .B(n817), .ZN(n911) );
  XNOR2_X1 U905 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NOR2_X1 U906 ( .A1(n911), .A2(n827), .ZN(n949) );
  NAND2_X1 U907 ( .A1(n949), .A2(n830), .ZN(n825) );
  NAND2_X1 U908 ( .A1(n818), .A2(n825), .ZN(n819) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n988) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n891), .ZN(n936) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n888), .ZN(n932) );
  NOR2_X1 U913 ( .A1(n820), .A2(n932), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U915 ( .A1(n936), .A2(n823), .ZN(n824) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n824), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n911), .A2(n827), .ZN(n947) );
  NAND2_X1 U919 ( .A1(n828), .A2(n947), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U921 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n834) );
  XNOR2_X1 U924 ( .A(KEYINPUT105), .B(n834), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n835), .A2(G661), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U928 ( .A(n838), .ZN(G319) );
  XNOR2_X1 U929 ( .A(G2427), .B(G1348), .ZN(n848) );
  XOR2_X1 U930 ( .A(G2451), .B(G2430), .Z(n840) );
  XNOR2_X1 U931 ( .A(G1341), .B(G2443), .ZN(n839) );
  XNOR2_X1 U932 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U933 ( .A(G2438), .B(G2435), .Z(n842) );
  XNOR2_X1 U934 ( .A(KEYINPUT103), .B(G2454), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U936 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U937 ( .A(KEYINPUT102), .B(G2446), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U939 ( .A(n848), .B(n847), .ZN(n849) );
  NAND2_X1 U940 ( .A1(n849), .A2(G14), .ZN(n850) );
  XOR2_X1 U941 ( .A(KEYINPUT104), .B(n850), .Z(G401) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n852) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U945 ( .A(G2678), .B(KEYINPUT42), .Z(n854) );
  XNOR2_X1 U946 ( .A(G2072), .B(KEYINPUT43), .ZN(n853) );
  XNOR2_X1 U947 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U948 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U950 ( .A(n858), .B(n857), .ZN(G227) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(KEYINPUT109), .Z(n860) );
  XNOR2_X1 U952 ( .A(G1961), .B(G1956), .ZN(n859) );
  XNOR2_X1 U953 ( .A(n860), .B(n859), .ZN(n870) );
  XOR2_X1 U954 ( .A(KEYINPUT110), .B(KEYINPUT108), .Z(n862) );
  XNOR2_X1 U955 ( .A(G1991), .B(G1986), .ZN(n861) );
  XNOR2_X1 U956 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U957 ( .A(G1976), .B(G1966), .Z(n864) );
  XNOR2_X1 U958 ( .A(G1981), .B(G1971), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U960 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U961 ( .A(G1996), .B(G2474), .ZN(n867) );
  XNOR2_X1 U962 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G124), .A2(n900), .ZN(n871) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(n871), .Z(n872) );
  XNOR2_X1 U966 ( .A(n872), .B(KEYINPUT111), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G100), .A2(n622), .ZN(n873) );
  NAND2_X1 U968 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U969 ( .A1(G112), .A2(n901), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G136), .A2(n905), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U972 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G130), .A2(n900), .ZN(n880) );
  NAND2_X1 U974 ( .A1(G118), .A2(n901), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U976 ( .A(KEYINPUT112), .B(n881), .ZN(n887) );
  NAND2_X1 U977 ( .A1(n622), .A2(G106), .ZN(n882) );
  XOR2_X1 U978 ( .A(KEYINPUT113), .B(n882), .Z(n884) );
  NAND2_X1 U979 ( .A1(n905), .A2(G142), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U981 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n899) );
  XOR2_X1 U984 ( .A(G164), .B(n930), .Z(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U986 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n893) );
  XNOR2_X1 U987 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U990 ( .A(G160), .B(G162), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n913) );
  NAND2_X1 U993 ( .A1(G127), .A2(n900), .ZN(n903) );
  NAND2_X1 U994 ( .A1(G115), .A2(n901), .ZN(n902) );
  NAND2_X1 U995 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U996 ( .A(n904), .B(KEYINPUT47), .ZN(n907) );
  NAND2_X1 U997 ( .A1(G139), .A2(n905), .ZN(n906) );
  NAND2_X1 U998 ( .A1(n907), .A2(n906), .ZN(n910) );
  NAND2_X1 U999 ( .A1(n622), .A2(G103), .ZN(n908) );
  XOR2_X1 U1000 ( .A(KEYINPUT114), .B(n908), .Z(n909) );
  NOR2_X1 U1001 ( .A1(n910), .A2(n909), .ZN(n939) );
  XNOR2_X1 U1002 ( .A(n911), .B(n939), .ZN(n912) );
  XNOR2_X1 U1003 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1005 ( .A(n986), .B(n915), .ZN(n917) );
  XNOR2_X1 U1006 ( .A(G286), .B(G171), .ZN(n916) );
  XNOR2_X1 U1007 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1008 ( .A(n918), .B(n980), .ZN(n919) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n919), .ZN(n920) );
  XOR2_X1 U1010 ( .A(KEYINPUT117), .B(n920), .Z(G397) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n922), .ZN(n923) );
  AND2_X1 U1014 ( .A1(G319), .A2(n923), .ZN(n925) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1016 ( .A1(n925), .A2(n924), .ZN(G225) );
  XOR2_X1 U1017 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  NOR2_X1 U1019 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1020 ( .A(n928), .B(KEYINPUT106), .ZN(G325) );
  XNOR2_X1 U1021 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U1022 ( .A(KEYINPUT55), .ZN(n976) );
  XOR2_X1 U1023 ( .A(G2084), .B(G160), .Z(n929) );
  NOR2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n934) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n946) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1029 ( .A(KEYINPUT119), .B(n937), .Z(n938) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n938), .Z(n944) );
  XOR2_X1 U1031 ( .A(G2072), .B(n939), .Z(n941) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(KEYINPUT50), .B(n942), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n951) );
  INV_X1 U1037 ( .A(n947), .ZN(n948) );
  NOR2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1039 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(KEYINPUT120), .B(n952), .ZN(n953) );
  XOR2_X1 U1041 ( .A(KEYINPUT52), .B(n953), .Z(n954) );
  NAND2_X1 U1042 ( .A1(n976), .A2(n954), .ZN(n955) );
  NAND2_X1 U1043 ( .A1(n955), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n971) );
  XOR2_X1 U1045 ( .A(G1991), .B(G25), .Z(n956) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(n956), .ZN(n968) );
  XNOR2_X1 U1047 ( .A(G27), .B(n957), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(G2067), .B(KEYINPUT122), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G26), .B(n958), .ZN(n959) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1054 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(KEYINPUT123), .B(n965), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(n966), .A2(G28), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(KEYINPUT53), .B(n969), .ZN(n970) );
  NOR2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1060 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1061 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1062 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1063 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1064 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1065 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n979), .ZN(n1033) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n1005) );
  XNOR2_X1 U1068 ( .A(n980), .B(G1341), .ZN(n985) );
  XOR2_X1 U1069 ( .A(G168), .B(G1966), .Z(n981) );
  NOR2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(KEYINPUT57), .B(n983), .ZN(n984) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n1003) );
  XNOR2_X1 U1073 ( .A(G1348), .B(n986), .ZN(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n995) );
  INV_X1 U1075 ( .A(G1971), .ZN(n989) );
  NOR2_X1 U1076 ( .A1(G166), .A2(n989), .ZN(n993) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n1000) );
  XNOR2_X1 U1080 ( .A(n996), .B(G1956), .ZN(n998) );
  XNOR2_X1 U1081 ( .A(G171), .B(G1961), .ZN(n997) );
  NAND2_X1 U1082 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1083 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(n1001), .B(KEYINPUT124), .ZN(n1002) );
  NAND2_X1 U1085 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1086 ( .A1(n1005), .A2(n1004), .ZN(n1031) );
  INV_X1 U1087 ( .A(G16), .ZN(n1029) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1090 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1091 ( .A(KEYINPUT126), .B(n1008), .Z(n1010) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1009) );
  NOR2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1011), .ZN(n1015) );
  XNOR2_X1 U1095 ( .A(G1961), .B(G5), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1012) );
  NOR2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1098 ( .A1(n1015), .A2(n1014), .ZN(n1026) );
  XNOR2_X1 U1099 ( .A(G1956), .B(G20), .ZN(n1020) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G6), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G19), .B(G1341), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XNOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(G4), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1112 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1113 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1114 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  XNOR2_X1 U1116 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1117 ( .A(G120), .ZN(G236) );
  INV_X1 U1118 ( .A(G96), .ZN(G221) );
  INV_X1 U1119 ( .A(G69), .ZN(G235) );
  INV_X1 U1120 ( .A(G171), .ZN(G301) );
  INV_X1 U1121 ( .A(G108), .ZN(G238) );
endmodule

