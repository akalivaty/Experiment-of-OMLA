

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782;

  XNOR2_X1 U368 ( .A(n569), .B(KEYINPUT31), .ZN(n702) );
  AND2_X1 U369 ( .A1(n741), .A2(n597), .ZN(n593) );
  INV_X1 U370 ( .A(n541), .ZN(n552) );
  AND2_X1 U371 ( .A1(n698), .A2(n603), .ZN(n605) );
  XNOR2_X1 U372 ( .A(n478), .B(n477), .ZN(n558) );
  OR2_X1 U373 ( .A1(n750), .A2(G902), .ZN(n398) );
  XNOR2_X1 U374 ( .A(n417), .B(n510), .ZN(n523) );
  XNOR2_X1 U375 ( .A(n451), .B(KEYINPUT80), .ZN(n453) );
  XNOR2_X1 U376 ( .A(G143), .B(G128), .ZN(n452) );
  XNOR2_X1 U377 ( .A(G125), .B(G140), .ZN(n404) );
  INV_X1 U378 ( .A(G953), .ZN(n771) );
  AND2_X2 U379 ( .A1(n444), .A2(KEYINPUT84), .ZN(n370) );
  OR2_X2 U380 ( .A1(n740), .A2(n423), .ZN(n418) );
  XNOR2_X2 U381 ( .A(n348), .B(n548), .ZN(n776) );
  NAND2_X1 U382 ( .A1(n420), .A2(n421), .ZN(n348) );
  INV_X2 U383 ( .A(KEYINPUT64), .ZN(n451) );
  NAND2_X1 U384 ( .A1(n349), .A2(n619), .ZN(n620) );
  NOR2_X2 U385 ( .A1(n617), .A2(n616), .ZN(n349) );
  NOR2_X1 U386 ( .A1(n667), .A2(n782), .ZN(n594) );
  BUF_X1 U387 ( .A(n566), .Z(n726) );
  XNOR2_X1 U388 ( .A(n593), .B(KEYINPUT42), .ZN(n782) );
  XNOR2_X2 U389 ( .A(n586), .B(KEYINPUT115), .ZN(n712) );
  INV_X2 U390 ( .A(n724), .ZN(n590) );
  XNOR2_X2 U391 ( .A(n398), .B(n362), .ZN(n724) );
  NOR2_X2 U392 ( .A1(n673), .A2(G902), .ZN(n415) );
  XNOR2_X2 U393 ( .A(n415), .B(G472), .ZN(n566) );
  XNOR2_X2 U394 ( .A(n592), .B(KEYINPUT1), .ZN(n541) );
  BUF_X2 U395 ( .A(n541), .Z(n720) );
  XNOR2_X2 U396 ( .A(n546), .B(KEYINPUT33), .ZN(n740) );
  NAND2_X2 U397 ( .A1(n552), .A2(n545), .ZN(n546) );
  INV_X4 U398 ( .A(G104), .ZN(n396) );
  INV_X1 U399 ( .A(n352), .ZN(n604) );
  INV_X1 U400 ( .A(KEYINPUT6), .ZN(n353) );
  INV_X1 U401 ( .A(KEYINPUT68), .ZN(n395) );
  XNOR2_X2 U402 ( .A(G107), .B(KEYINPUT73), .ZN(n405) );
  AND2_X1 U403 ( .A1(n374), .A2(n372), .ZN(n371) );
  NAND2_X1 U404 ( .A1(n445), .A2(n370), .ZN(n369) );
  XNOR2_X1 U405 ( .A(n385), .B(n585), .ZN(n667) );
  NOR2_X1 U406 ( .A1(n778), .A2(n695), .ZN(n614) );
  XNOR2_X1 U407 ( .A(n354), .B(KEYINPUT116), .ZN(n778) );
  NAND2_X1 U408 ( .A1(n382), .A2(n379), .ZN(n632) );
  XNOR2_X1 U409 ( .A(n599), .B(n598), .ZN(n692) );
  NAND2_X1 U410 ( .A1(n577), .A2(n576), .ZN(n583) );
  XNOR2_X1 U411 ( .A(n428), .B(n559), .ZN(n703) );
  XNOR2_X1 U412 ( .A(n523), .B(KEYINPUT95), .ZN(n766) );
  XNOR2_X1 U413 ( .A(n492), .B(n491), .ZN(n521) );
  XNOR2_X1 U414 ( .A(n488), .B(n394), .ZN(n434) );
  XNOR2_X1 U415 ( .A(n395), .B(KEYINPUT16), .ZN(n394) );
  XNOR2_X1 U416 ( .A(n405), .B(G110), .ZN(n511) );
  XNOR2_X1 U417 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n483) );
  XOR2_X1 U418 ( .A(KEYINPUT92), .B(KEYINPUT18), .Z(n484) );
  XNOR2_X2 U419 ( .A(n350), .B(G469), .ZN(n592) );
  NOR2_X1 U420 ( .A1(n680), .A2(G902), .ZN(n350) );
  BUF_X1 U421 ( .A(n709), .Z(n351) );
  XNOR2_X1 U422 ( .A(n608), .B(n584), .ZN(n709) );
  XNOR2_X1 U423 ( .A(n566), .B(n353), .ZN(n352) );
  AND2_X1 U424 ( .A1(n401), .A2(n552), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n435), .B(KEYINPUT111), .ZN(n355) );
  XNOR2_X1 U426 ( .A(n482), .B(n481), .ZN(n356) );
  XNOR2_X1 U427 ( .A(n482), .B(n481), .ZN(n417) );
  XNOR2_X1 U428 ( .A(n387), .B(KEYINPUT45), .ZN(n648) );
  NOR2_X2 U429 ( .A1(n671), .A2(n754), .ZN(n672) );
  NOR2_X2 U430 ( .A1(n649), .A2(n409), .ZN(n706) );
  NOR2_X2 U431 ( .A1(n676), .A2(n754), .ZN(n678) );
  NOR2_X2 U432 ( .A1(n664), .A2(n754), .ZN(n665) );
  NOR2_X2 U433 ( .A1(n655), .A2(n754), .ZN(n657) );
  NOR2_X1 U434 ( .A1(n720), .A2(n567), .ZN(n450) );
  XNOR2_X2 U435 ( .A(n497), .B(n496), .ZN(n608) );
  NAND2_X1 U436 ( .A1(n355), .A2(n570), .ZN(n393) );
  XNOR2_X1 U437 ( .A(n479), .B(n386), .ZN(n723) );
  XNOR2_X1 U438 ( .A(KEYINPUT101), .B(KEYINPUT21), .ZN(n386) );
  XNOR2_X1 U439 ( .A(n620), .B(n367), .ZN(n449) );
  XNOR2_X1 U440 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  INV_X1 U441 ( .A(KEYINPUT85), .ZN(n448) );
  INV_X1 U442 ( .A(G237), .ZN(n493) );
  XOR2_X1 U443 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n455) );
  XNOR2_X1 U444 ( .A(G116), .B(G107), .ZN(n457) );
  XOR2_X1 U445 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n458) );
  NOR2_X1 U446 ( .A1(G953), .A2(G237), .ZN(n517) );
  XNOR2_X1 U447 ( .A(n404), .B(n403), .ZN(n765) );
  INV_X1 U448 ( .A(KEYINPUT10), .ZN(n403) );
  INV_X1 U449 ( .A(G137), .ZN(n507) );
  INV_X1 U450 ( .A(n377), .ZN(n445) );
  NAND2_X1 U451 ( .A1(n389), .A2(n361), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n391) );
  NAND2_X1 U453 ( .A1(n590), .A2(n589), .ZN(n397) );
  XOR2_X1 U454 ( .A(KEYINPUT3), .B(G119), .Z(n491) );
  XNOR2_X1 U455 ( .A(G137), .B(G128), .ZN(n524) );
  XNOR2_X1 U456 ( .A(n765), .B(G146), .ZN(n533) );
  NAND2_X1 U457 ( .A1(n381), .A2(n380), .ZN(n379) );
  AND2_X1 U458 ( .A1(n384), .A2(n383), .ZN(n382) );
  NOR2_X1 U459 ( .A1(n622), .A2(n606), .ZN(n402) );
  BUF_X1 U460 ( .A(n561), .Z(n568) );
  XNOR2_X1 U461 ( .A(n476), .B(G475), .ZN(n477) );
  NOR2_X1 U462 ( .A1(n668), .A2(G902), .ZN(n478) );
  XNOR2_X1 U463 ( .A(n464), .B(n463), .ZN(n556) );
  INV_X1 U464 ( .A(KEYINPUT47), .ZN(n426) );
  XNOR2_X1 U465 ( .A(n368), .B(KEYINPUT20), .ZN(n534) );
  AND2_X1 U466 ( .A1(n447), .A2(n658), .ZN(n446) );
  NAND2_X1 U467 ( .A1(n777), .A2(n448), .ZN(n447) );
  INV_X1 U468 ( .A(KEYINPUT88), .ZN(n392) );
  XNOR2_X1 U469 ( .A(n571), .B(n390), .ZN(n389) );
  INV_X1 U470 ( .A(KEYINPUT89), .ZN(n390) );
  XNOR2_X1 U471 ( .A(n495), .B(KEYINPUT81), .ZN(n496) );
  XNOR2_X1 U472 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n526) );
  INV_X1 U473 ( .A(KEYINPUT67), .ZN(n466) );
  XOR2_X1 U474 ( .A(G125), .B(KEYINPUT17), .Z(n486) );
  XNOR2_X1 U475 ( .A(KEYINPUT4), .B(G146), .ZN(n481) );
  NAND2_X1 U476 ( .A1(G234), .A2(G237), .ZN(n500) );
  AND2_X1 U477 ( .A1(n633), .A2(n448), .ZN(n373) );
  NAND2_X1 U478 ( .A1(n498), .A2(G214), .ZN(n708) );
  NOR2_X1 U479 ( .A1(n583), .A2(n366), .ZN(n380) );
  INV_X1 U480 ( .A(G902), .ZN(n494) );
  XOR2_X1 U481 ( .A(G134), .B(G122), .Z(n459) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n470) );
  XNOR2_X1 U483 ( .A(n465), .B(G113), .ZN(n425) );
  INV_X1 U484 ( .A(KEYINPUT28), .ZN(n407) );
  NOR2_X1 U485 ( .A1(n583), .A2(n582), .ZN(n607) );
  INV_X1 U486 ( .A(KEYINPUT22), .ZN(n441) );
  AND2_X1 U487 ( .A1(n711), .A2(n363), .ZN(n443) );
  XNOR2_X1 U488 ( .A(n532), .B(n530), .ZN(n399) );
  XNOR2_X1 U489 ( .A(G119), .B(G110), .ZN(n530) );
  NAND2_X1 U490 ( .A1(n378), .A2(n698), .ZN(n385) );
  INV_X1 U491 ( .A(n632), .ZN(n378) );
  INV_X1 U492 ( .A(KEYINPUT35), .ZN(n548) );
  NOR2_X1 U493 ( .A1(n422), .A2(n357), .ZN(n421) );
  NAND2_X1 U494 ( .A1(n556), .A2(n429), .ZN(n428) );
  INV_X1 U495 ( .A(n558), .ZN(n429) );
  OR2_X1 U496 ( .A1(n703), .A2(n698), .ZN(n427) );
  XOR2_X1 U497 ( .A(KEYINPUT77), .B(n611), .Z(n357) );
  XOR2_X1 U498 ( .A(n529), .B(n528), .Z(n358) );
  XOR2_X1 U499 ( .A(n484), .B(n483), .Z(n359) );
  AND2_X1 U500 ( .A1(n630), .A2(KEYINPUT85), .ZN(n360) );
  AND2_X1 U501 ( .A1(n572), .A2(n776), .ZN(n361) );
  XOR2_X1 U502 ( .A(n536), .B(n535), .Z(n362) );
  XOR2_X1 U503 ( .A(n723), .B(n480), .Z(n363) );
  AND2_X1 U504 ( .A1(n427), .A2(n426), .ZN(n364) );
  INV_X1 U505 ( .A(n777), .ZN(n630) );
  XNOR2_X1 U506 ( .A(n629), .B(n628), .ZN(n777) );
  NAND2_X1 U507 ( .A1(n568), .A2(n547), .ZN(n365) );
  XNOR2_X1 U508 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n366) );
  INV_X1 U509 ( .A(n547), .ZN(n423) );
  XOR2_X1 U510 ( .A(KEYINPUT86), .B(KEYINPUT48), .Z(n367) );
  NAND2_X1 U511 ( .A1(n641), .A2(G234), .ZN(n368) );
  NAND2_X1 U512 ( .A1(n371), .A2(n369), .ZN(n767) );
  NAND2_X1 U513 ( .A1(n376), .A2(n448), .ZN(n444) );
  NAND2_X1 U514 ( .A1(n376), .A2(n373), .ZN(n372) );
  NAND2_X1 U515 ( .A1(n377), .A2(n633), .ZN(n374) );
  NAND2_X1 U516 ( .A1(n375), .A2(n446), .ZN(n377) );
  NAND2_X1 U517 ( .A1(n449), .A2(n360), .ZN(n375) );
  INV_X1 U518 ( .A(n449), .ZN(n376) );
  INV_X1 U519 ( .A(n411), .ZN(n381) );
  NAND2_X1 U520 ( .A1(n583), .A2(n366), .ZN(n383) );
  NAND2_X1 U521 ( .A1(n411), .A2(n366), .ZN(n384) );
  NAND2_X1 U522 ( .A1(n391), .A2(n388), .ZN(n387) );
  XNOR2_X2 U523 ( .A(n396), .B(G122), .ZN(n488) );
  INV_X1 U524 ( .A(n397), .ZN(n603) );
  NOR2_X1 U525 ( .A1(n726), .A2(n397), .ZN(n408) );
  XNOR2_X1 U526 ( .A(n400), .B(n399), .ZN(n750) );
  XNOR2_X1 U527 ( .A(n358), .B(n533), .ZN(n400) );
  XNOR2_X1 U528 ( .A(n402), .B(KEYINPUT36), .ZN(n401) );
  BUF_X1 U529 ( .A(n595), .Z(n406) );
  XNOR2_X1 U530 ( .A(n408), .B(n407), .ZN(n591) );
  NAND2_X1 U531 ( .A1(n445), .A2(n444), .ZN(n409) );
  INV_X1 U532 ( .A(n582), .ZN(n410) );
  NAND2_X1 U533 ( .A1(n351), .A2(n410), .ZN(n411) );
  NAND2_X1 U534 ( .A1(n419), .A2(n418), .ZN(n420) );
  NOR2_X1 U535 ( .A1(n650), .A2(n706), .ZN(n412) );
  NOR2_X2 U536 ( .A1(n650), .A2(n706), .ZN(n413) );
  BUF_X1 U537 ( .A(n724), .Z(n414) );
  NOR2_X2 U538 ( .A1(n551), .A2(n538), .ZN(n539) );
  XNOR2_X1 U539 ( .A(n587), .B(KEYINPUT41), .ZN(n741) );
  NAND2_X1 U540 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X1 U541 ( .A(n409), .B(n633), .ZN(n416) );
  XNOR2_X1 U542 ( .A(n760), .B(n433), .ZN(n659) );
  XNOR2_X1 U543 ( .A(n430), .B(n356), .ZN(n433) );
  NAND2_X1 U544 ( .A1(n365), .A2(n740), .ZN(n419) );
  NOR2_X1 U545 ( .A1(n568), .A2(n547), .ZN(n422) );
  INV_X1 U546 ( .A(n488), .ZN(n424) );
  XNOR2_X1 U547 ( .A(n359), .B(n487), .ZN(n430) );
  XNOR2_X2 U548 ( .A(n431), .B(n521), .ZN(n760) );
  XNOR2_X2 U549 ( .A(n434), .B(n432), .ZN(n431) );
  INV_X1 U550 ( .A(n511), .ZN(n432) );
  INV_X1 U551 ( .A(n684), .ZN(n436) );
  NAND2_X1 U552 ( .A1(n438), .A2(n427), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n440), .A2(n439), .ZN(n438) );
  INV_X1 U554 ( .A(n702), .ZN(n439) );
  INV_X1 U555 ( .A(n685), .ZN(n440) );
  INV_X1 U556 ( .A(n554), .ZN(n551) );
  XNOR2_X2 U557 ( .A(n442), .B(n441), .ZN(n554) );
  NAND2_X1 U558 ( .A1(n561), .A2(n443), .ZN(n442) );
  NAND2_X1 U559 ( .A1(n705), .A2(n638), .ZN(n645) );
  NOR2_X1 U560 ( .A1(n705), .A2(KEYINPUT82), .ZN(n647) );
  AND2_X2 U561 ( .A1(n767), .A2(n648), .ZN(n705) );
  AND2_X2 U562 ( .A1(n558), .A2(n557), .ZN(n698) );
  BUF_X1 U563 ( .A(n685), .Z(n687) );
  NOR2_X1 U564 ( .A1(n592), .A2(n591), .ZN(n597) );
  XNOR2_X1 U565 ( .A(n470), .B(n469), .ZN(n475) );
  INV_X1 U566 ( .A(KEYINPUT105), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n468), .B(n467), .ZN(n469) );
  AND2_X1 U568 ( .A1(n597), .A2(n596), .ZN(n599) );
  BUF_X1 U569 ( .A(n412), .Z(n749) );
  BUF_X1 U570 ( .A(n692), .Z(n696) );
  INV_X1 U571 ( .A(KEYINPUT123), .ZN(n656) );
  XNOR2_X1 U572 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n540) );
  XNOR2_X2 U573 ( .A(n453), .B(n452), .ZN(n482) );
  NAND2_X1 U574 ( .A1(G234), .A2(n771), .ZN(n454) );
  XNOR2_X1 U575 ( .A(n455), .B(n454), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G217), .A2(n531), .ZN(n456) );
  XNOR2_X1 U577 ( .A(n482), .B(n456), .ZN(n462) );
  XNOR2_X1 U578 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U579 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U580 ( .A(n462), .B(n461), .ZN(n651) );
  NAND2_X1 U581 ( .A1(n651), .A2(n494), .ZN(n464) );
  XOR2_X1 U582 ( .A(KEYINPUT109), .B(G478), .Z(n463) );
  NAND2_X1 U583 ( .A1(G214), .A2(n517), .ZN(n465) );
  XNOR2_X1 U584 ( .A(n466), .B(G131), .ZN(n509) );
  XNOR2_X1 U585 ( .A(n509), .B(G143), .ZN(n468) );
  XOR2_X1 U586 ( .A(KEYINPUT106), .B(KEYINPUT11), .Z(n472) );
  XNOR2_X1 U587 ( .A(KEYINPUT107), .B(KEYINPUT12), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U589 ( .A(n533), .B(n473), .ZN(n474) );
  XNOR2_X1 U590 ( .A(n475), .B(n474), .ZN(n668) );
  XNOR2_X1 U591 ( .A(KEYINPUT13), .B(KEYINPUT108), .ZN(n476) );
  NOR2_X1 U592 ( .A1(n556), .A2(n558), .ZN(n711) );
  NAND2_X1 U593 ( .A1(n534), .A2(G221), .ZN(n479) );
  INV_X1 U594 ( .A(KEYINPUT102), .ZN(n480) );
  NAND2_X1 U595 ( .A1(G224), .A2(n771), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U597 ( .A(KEYINPUT91), .B(G101), .ZN(n490) );
  XNOR2_X1 U598 ( .A(G116), .B(G113), .ZN(n489) );
  XNOR2_X1 U599 ( .A(n490), .B(n489), .ZN(n492) );
  NAND2_X1 U600 ( .A1(n659), .A2(n641), .ZN(n497) );
  NAND2_X1 U601 ( .A1(n494), .A2(n493), .ZN(n498) );
  NAND2_X1 U602 ( .A1(n498), .A2(G210), .ZN(n495) );
  NAND2_X1 U603 ( .A1(n608), .A2(n708), .ZN(n606) );
  XOR2_X1 U604 ( .A(KEYINPUT74), .B(KEYINPUT19), .Z(n499) );
  XNOR2_X1 U605 ( .A(n606), .B(n499), .ZN(n595) );
  XNOR2_X1 U606 ( .A(n500), .B(KEYINPUT14), .ZN(n501) );
  NAND2_X1 U607 ( .A1(G952), .A2(n501), .ZN(n739) );
  NOR2_X1 U608 ( .A1(n739), .A2(G953), .ZN(n580) );
  AND2_X1 U609 ( .A1(G902), .A2(n501), .ZN(n578) );
  NOR2_X1 U610 ( .A1(G898), .A2(n771), .ZN(n762) );
  NAND2_X1 U611 ( .A1(n578), .A2(n762), .ZN(n502) );
  XNOR2_X1 U612 ( .A(KEYINPUT93), .B(n502), .ZN(n503) );
  NOR2_X1 U613 ( .A1(n580), .A2(n503), .ZN(n504) );
  XNOR2_X1 U614 ( .A(n504), .B(KEYINPUT94), .ZN(n505) );
  NOR2_X2 U615 ( .A1(n595), .A2(n505), .ZN(n506) );
  XNOR2_X2 U616 ( .A(n506), .B(KEYINPUT0), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n507), .B(G134), .ZN(n508) );
  XNOR2_X1 U618 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U619 ( .A(G101), .B(n511), .Z(n515) );
  NAND2_X1 U620 ( .A1(G227), .A2(n771), .ZN(n512) );
  XNOR2_X1 U621 ( .A(G140), .B(n512), .ZN(n513) );
  XNOR2_X1 U622 ( .A(n513), .B(G104), .ZN(n514) );
  XNOR2_X1 U623 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U624 ( .A(n766), .B(n516), .ZN(n680) );
  XNOR2_X1 U625 ( .A(KEYINPUT72), .B(KEYINPUT5), .ZN(n519) );
  NAND2_X1 U626 ( .A1(G210), .A2(n517), .ZN(n518) );
  XNOR2_X1 U627 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U628 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U629 ( .A(n523), .B(n522), .ZN(n673) );
  XOR2_X1 U630 ( .A(KEYINPUT24), .B(KEYINPUT96), .Z(n525) );
  XNOR2_X1 U631 ( .A(n525), .B(n524), .ZN(n529) );
  XOR2_X1 U632 ( .A(KEYINPUT98), .B(KEYINPUT23), .Z(n527) );
  XNOR2_X1 U633 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U634 ( .A1(G221), .A2(n531), .ZN(n532) );
  NAND2_X1 U635 ( .A1(n534), .A2(G217), .ZN(n536) );
  XNOR2_X1 U636 ( .A(KEYINPUT25), .B(KEYINPUT100), .ZN(n535) );
  NOR2_X1 U637 ( .A1(n604), .A2(n414), .ZN(n537) );
  NAND2_X1 U638 ( .A1(n552), .A2(n537), .ZN(n538) );
  XNOR2_X1 U639 ( .A(n540), .B(n539), .ZN(n780) );
  NAND2_X1 U640 ( .A1(n720), .A2(n726), .ZN(n542) );
  NOR2_X1 U641 ( .A1(n551), .A2(n542), .ZN(n543) );
  NAND2_X1 U642 ( .A1(n543), .A2(n590), .ZN(n691) );
  AND2_X1 U643 ( .A1(n780), .A2(n691), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n556), .A2(n558), .ZN(n611) );
  AND2_X1 U645 ( .A1(n724), .A2(n363), .ZN(n718) );
  INV_X1 U646 ( .A(n718), .ZN(n716) );
  INV_X1 U647 ( .A(n604), .ZN(n544) );
  NOR2_X1 U648 ( .A1(n716), .A2(n544), .ZN(n545) );
  XOR2_X1 U649 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n547) );
  NAND2_X1 U650 ( .A1(n571), .A2(n776), .ZN(n550) );
  NAND2_X1 U651 ( .A1(n550), .A2(KEYINPUT44), .ZN(n570) );
  NOR2_X1 U652 ( .A1(n552), .A2(n604), .ZN(n553) );
  NAND2_X1 U653 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U654 ( .A1(n590), .A2(n555), .ZN(n684) );
  INV_X1 U655 ( .A(n556), .ZN(n557) );
  INV_X1 U656 ( .A(KEYINPUT110), .ZN(n559) );
  NOR2_X1 U657 ( .A1(n716), .A2(n592), .ZN(n560) );
  NAND2_X1 U658 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U659 ( .A(n562), .B(KEYINPUT103), .ZN(n563) );
  NAND2_X1 U660 ( .A1(n563), .A2(n726), .ZN(n565) );
  INV_X1 U661 ( .A(KEYINPUT104), .ZN(n564) );
  XNOR2_X1 U662 ( .A(n565), .B(n564), .ZN(n685) );
  INV_X1 U663 ( .A(n566), .ZN(n573) );
  NAND2_X1 U664 ( .A1(n718), .A2(n573), .ZN(n567) );
  NAND2_X1 U665 ( .A1(n568), .A2(n450), .ZN(n569) );
  INV_X1 U666 ( .A(KEYINPUT44), .ZN(n572) );
  NAND2_X1 U667 ( .A1(n573), .A2(n708), .ZN(n575) );
  XNOR2_X1 U668 ( .A(KEYINPUT113), .B(KEYINPUT30), .ZN(n574) );
  XNOR2_X1 U669 ( .A(n575), .B(n574), .ZN(n577) );
  INV_X1 U670 ( .A(n592), .ZN(n576) );
  NAND2_X1 U671 ( .A1(G953), .A2(n578), .ZN(n579) );
  NOR2_X1 U672 ( .A1(n579), .A2(G900), .ZN(n581) );
  OR2_X1 U673 ( .A1(n581), .A2(n580), .ZN(n588) );
  NAND2_X1 U674 ( .A1(n718), .A2(n588), .ZN(n582) );
  XNOR2_X1 U675 ( .A(KEYINPUT71), .B(KEYINPUT38), .ZN(n584) );
  INV_X1 U676 ( .A(KEYINPUT40), .ZN(n585) );
  NAND2_X1 U677 ( .A1(n708), .A2(n709), .ZN(n586) );
  NAND2_X1 U678 ( .A1(n712), .A2(n711), .ZN(n587) );
  AND2_X1 U679 ( .A1(n723), .A2(n588), .ZN(n589) );
  XNOR2_X1 U680 ( .A(n594), .B(KEYINPUT46), .ZN(n619) );
  INV_X1 U681 ( .A(n406), .ZN(n596) );
  INV_X1 U682 ( .A(KEYINPUT79), .ZN(n598) );
  XNOR2_X1 U683 ( .A(KEYINPUT70), .B(n364), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n692), .A2(n600), .ZN(n601) );
  XNOR2_X1 U685 ( .A(n601), .B(KEYINPUT69), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n427), .A2(n692), .ZN(n602) );
  NAND2_X1 U687 ( .A1(KEYINPUT47), .A2(n602), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n622) );
  BUF_X1 U689 ( .A(n608), .Z(n626) );
  NAND2_X1 U690 ( .A1(n607), .A2(n626), .ZN(n610) );
  INV_X1 U691 ( .A(KEYINPUT114), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n610), .B(n609), .ZN(n613) );
  INV_X1 U693 ( .A(n611), .ZN(n612) );
  AND2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n695) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U696 ( .A(n708), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n623), .A2(n720), .ZN(n625) );
  INV_X1 U699 ( .A(KEYINPUT43), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(n627) );
  OR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n629) );
  INV_X1 U702 ( .A(KEYINPUT112), .ZN(n628) );
  INV_X1 U703 ( .A(n703), .ZN(n631) );
  OR2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n658) );
  INV_X1 U705 ( .A(KEYINPUT84), .ZN(n633) );
  INV_X1 U706 ( .A(n641), .ZN(n636) );
  NAND2_X1 U707 ( .A1(KEYINPUT2), .A2(KEYINPUT83), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n634), .A2(KEYINPUT82), .ZN(n635) );
  NOR2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n643) );
  INV_X1 U710 ( .A(n643), .ZN(n637) );
  AND2_X1 U711 ( .A1(KEYINPUT82), .A2(n637), .ZN(n638) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n639), .A2(KEYINPUT83), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  OR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U717 ( .A1(n646), .A2(n647), .ZN(n650) );
  BUF_X1 U718 ( .A(n648), .Z(n755) );
  NAND2_X1 U719 ( .A1(n755), .A2(KEYINPUT2), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n413), .A2(G478), .ZN(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT122), .B(n651), .Z(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n655) );
  INV_X1 U723 ( .A(G952), .ZN(n654) );
  AND2_X1 U724 ( .A1(n654), .A2(G953), .ZN(n754) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(G63) );
  XNOR2_X1 U726 ( .A(n658), .B(G134), .ZN(G36) );
  NAND2_X1 U727 ( .A1(n413), .A2(G210), .ZN(n663) );
  BUF_X1 U728 ( .A(n659), .Z(n661) );
  XNOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U733 ( .A(G131), .B(KEYINPUT127), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(G33) );
  NAND2_X1 U735 ( .A1(n412), .A2(G475), .ZN(n670) );
  XOR2_X1 U736 ( .A(KEYINPUT59), .B(n668), .Z(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U739 ( .A1(n413), .A2(G472), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n673), .B(KEYINPUT62), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U742 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n677) );
  XNOR2_X1 U743 ( .A(n678), .B(n677), .ZN(G57) );
  NAND2_X1 U744 ( .A1(n749), .A2(G469), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U748 ( .A1(n683), .A2(n754), .ZN(G54) );
  XOR2_X1 U749 ( .A(G101), .B(n684), .Z(G3) );
  NAND2_X1 U750 ( .A1(n687), .A2(n698), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(G104), .ZN(G6) );
  XOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U753 ( .A1(n687), .A2(n703), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U755 ( .A(G107), .B(n690), .ZN(G9) );
  XNOR2_X1 U756 ( .A(G110), .B(n691), .ZN(G12) );
  XOR2_X1 U757 ( .A(G128), .B(KEYINPUT29), .Z(n694) );
  NAND2_X1 U758 ( .A1(n696), .A2(n703), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n694), .B(n693), .ZN(G30) );
  XOR2_X1 U760 ( .A(G143), .B(n695), .Z(G45) );
  NAND2_X1 U761 ( .A1(n696), .A2(n698), .ZN(n697) );
  XNOR2_X1 U762 ( .A(n697), .B(G146), .ZN(G48) );
  XOR2_X1 U763 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n700) );
  NAND2_X1 U764 ( .A1(n702), .A2(n698), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(G113), .B(n701), .ZN(G15) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U768 ( .A(n704), .B(G116), .ZN(G18) );
  NOR2_X1 U769 ( .A1(n705), .A2(KEYINPUT2), .ZN(n707) );
  OR2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n746) );
  OR2_X1 U771 ( .A1(n351), .A2(n708), .ZN(n710) );
  NAND2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U773 ( .A1(n712), .A2(n427), .ZN(n713) );
  NAND2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U775 ( .A1(n715), .A2(n740), .ZN(n735) );
  NAND2_X1 U776 ( .A1(n720), .A2(n716), .ZN(n717) );
  NAND2_X1 U777 ( .A1(n717), .A2(KEYINPUT50), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n718), .A2(KEYINPUT50), .ZN(n719) );
  NAND2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n414), .A2(n723), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n725), .B(KEYINPUT49), .ZN(n727) );
  NAND2_X1 U783 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n730), .A2(n450), .ZN(n731) );
  XOR2_X1 U786 ( .A(KEYINPUT119), .B(n731), .Z(n732) );
  XNOR2_X1 U787 ( .A(KEYINPUT51), .B(n732), .ZN(n733) );
  NAND2_X1 U788 ( .A1(n733), .A2(n741), .ZN(n734) );
  NAND2_X1 U789 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n736), .B(KEYINPUT52), .ZN(n737) );
  XOR2_X1 U791 ( .A(KEYINPUT120), .B(n737), .Z(n738) );
  NOR2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n744) );
  AND2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U794 ( .A(KEYINPUT121), .B(n742), .Z(n743) );
  NOR2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U797 ( .A1(n747), .A2(G953), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n748), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U799 ( .A1(n749), .A2(G217), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n750), .B(KEYINPUT124), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U802 ( .A1(n754), .A2(n753), .ZN(G66) );
  NAND2_X1 U803 ( .A1(n771), .A2(n755), .ZN(n759) );
  NAND2_X1 U804 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U805 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n764) );
  XOR2_X1 U808 ( .A(n760), .B(KEYINPUT125), .Z(n761) );
  NOR2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U811 ( .A(n766), .B(n765), .ZN(n769) );
  XNOR2_X1 U812 ( .A(n416), .B(n769), .ZN(n768) );
  NOR2_X1 U813 ( .A1(n768), .A2(G953), .ZN(n774) );
  XOR2_X1 U814 ( .A(G227), .B(n769), .Z(n770) );
  NAND2_X1 U815 ( .A1(n770), .A2(G900), .ZN(n772) );
  NOR2_X1 U816 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U817 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U818 ( .A(KEYINPUT126), .B(n775), .ZN(G72) );
  XNOR2_X1 U819 ( .A(n776), .B(G122), .ZN(G24) );
  XOR2_X1 U820 ( .A(G140), .B(n777), .Z(G42) );
  XNOR2_X1 U821 ( .A(G125), .B(KEYINPUT37), .ZN(n779) );
  XNOR2_X1 U822 ( .A(n779), .B(n778), .ZN(G27) );
  BUF_X1 U823 ( .A(n780), .Z(n781) );
  XNOR2_X1 U824 ( .A(G119), .B(n781), .ZN(G21) );
  XOR2_X1 U825 ( .A(n782), .B(G137), .Z(G39) );
endmodule

