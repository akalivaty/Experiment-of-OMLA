//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT75), .A2(G125), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT75), .A2(G125), .ZN(new_n194));
  OAI21_X1  g008(.A(G140), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(G125), .A2(G140), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(new_n194), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n191), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT75), .B(G125), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n192), .A3(new_n200), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n196), .B1(new_n204), .B2(G140), .ZN(new_n206));
  OAI211_X1 g020(.A(G146), .B(new_n205), .C1(new_n206), .C2(new_n192), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(G128), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n210), .B(new_n212), .C1(new_n213), .C2(KEYINPUT23), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n214), .B2(new_n215), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT24), .B(G110), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT73), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(G119), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n212), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n212), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT73), .B1(new_n224), .B2(new_n219), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n216), .A2(new_n218), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n208), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  XNOR2_X1  g042(.A(G125), .B(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n191), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n214), .A2(G110), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n224), .A2(new_n219), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n207), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n227), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n228), .B1(new_n227), .B2(new_n233), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n190), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n190), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n227), .A2(new_n233), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(KEYINPUT76), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(G234), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G902), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n242), .A3(new_n239), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n242), .A4(new_n239), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n248), .A2(KEYINPUT77), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT77), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n251), .A3(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n243), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n245), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G472), .A2(G902), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n255), .B(KEYINPUT71), .Z(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT65), .B1(new_n258), .B2(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n191), .A3(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(G146), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT0), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(new_n209), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT64), .B1(new_n264), .B2(new_n209), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n263), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n263), .B2(new_n267), .ZN(new_n271));
  INV_X1    g085(.A(new_n265), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(G137), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  INV_X1    g096(.A(G131), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n279), .A3(new_n283), .A4(new_n280), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(KEYINPUT66), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n286), .A3(G131), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(KEYINPUT68), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT68), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n274), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n191), .A2(G143), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n262), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n270), .A2(new_n295), .A3(new_n291), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n263), .B1(new_n298), .B2(new_n209), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n280), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n276), .A2(G137), .ZN(new_n302));
  OAI21_X1  g116(.A(G131), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(new_n284), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G113), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT2), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G113), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n211), .A2(G116), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n307), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n309), .ZN(new_n314));
  XNOR2_X1  g128(.A(G116), .B(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n305), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT28), .B1(new_n290), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n285), .A2(new_n287), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n305), .B1(new_n273), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n317), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n285), .A2(KEYINPUT68), .A3(new_n287), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n273), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n321), .B1(new_n329), .B2(KEYINPUT28), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G210), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT27), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G101), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n257), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n335), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n290), .A2(new_n320), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n324), .ZN(new_n340));
  OAI211_X1 g154(.A(KEYINPUT70), .B(new_n337), .C1(new_n340), .C2(new_n321), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n323), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n317), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n300), .B2(new_n304), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT69), .B1(new_n328), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n290), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n346), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n335), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n343), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n318), .B1(new_n323), .B2(new_n344), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n290), .A2(new_n350), .A3(new_n347), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n350), .B1(new_n290), .B2(new_n347), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n353), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT31), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n256), .B1(new_n342), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n336), .A2(new_n341), .B1(new_n354), .B2(new_n360), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT32), .B1(new_n365), .B2(new_n256), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n339), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n349), .A2(new_n351), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n355), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT72), .B1(new_n370), .B2(new_n335), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n358), .A2(new_n339), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT72), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n337), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT29), .B1(new_n330), .B2(new_n335), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n300), .A2(new_n304), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n317), .B1(new_n328), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n339), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n321), .B1(new_n379), .B2(KEYINPUT28), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n335), .A2(KEYINPUT29), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G472), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n254), .B1(new_n367), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G475), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n188), .A3(G214), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n258), .ZN(new_n389));
  AOI21_X1  g203(.A(G143), .B1(new_n331), .B2(G214), .ZN(new_n390));
  OAI21_X1  g204(.A(G131), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n258), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n331), .A2(G143), .A3(G214), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n283), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n394), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT17), .A3(G131), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n203), .A2(new_n396), .A3(new_n207), .A4(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(G104), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n195), .A2(new_n197), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n230), .B1(new_n403), .B2(new_n191), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n393), .A2(new_n394), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(KEYINPUT18), .A3(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n399), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n402), .B1(new_n399), .B2(new_n408), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n386), .B1(new_n411), .B2(new_n242), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n391), .A2(new_n395), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n195), .A2(KEYINPUT19), .A3(new_n197), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT19), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n229), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n191), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n207), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n408), .ZN(new_n419));
  INV_X1    g233(.A(new_n402), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n399), .A2(new_n402), .A3(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n422), .A3(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT20), .ZN(new_n429));
  NOR3_X1   g243(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n421), .B2(new_n422), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT88), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n412), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT92), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n242), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G952), .ZN(new_n440));
  AOI211_X1 g254(.A(G953), .B(new_n440), .C1(G234), .C2(G237), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n310), .A2(G122), .ZN(new_n447));
  INV_X1    g261(.A(G107), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n258), .A2(G128), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n209), .A2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G134), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n276), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n446), .B1(new_n447), .B2(KEYINPUT14), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n445), .A2(G116), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n447), .A2(KEYINPUT89), .A3(KEYINPUT14), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n449), .B(new_n455), .C1(new_n462), .C2(new_n448), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT13), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n209), .B2(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n451), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n450), .A2(new_n464), .ZN(new_n467));
  OAI21_X1  g281(.A(G134), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n310), .A2(G122), .ZN(new_n469));
  OAI21_X1  g283(.A(G107), .B1(new_n469), .B2(new_n458), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n449), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n471), .A3(new_n454), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n241), .A3(G953), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n463), .B2(new_n472), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n444), .B(new_n242), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n479));
  NOR2_X1   g293(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n480));
  OAI21_X1  g294(.A(G478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n478), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n434), .A2(new_n443), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT78), .ZN(new_n486));
  INV_X1    g300(.A(G469), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n242), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n489));
  INV_X1    g303(.A(new_n270), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(KEYINPUT1), .C1(new_n258), .C2(G146), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G128), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n292), .B2(KEYINPUT1), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n297), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n448), .A2(G104), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n401), .A2(G107), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT3), .B1(new_n401), .B2(G107), .ZN(new_n501));
  AOI21_X1  g315(.A(G101), .B1(new_n401), .B2(G107), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT3), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n448), .A3(G104), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n502), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n500), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT82), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n496), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n496), .B2(new_n509), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n489), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n288), .A2(new_n289), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n501), .A2(new_n504), .A3(new_n499), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(G101), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n506), .A2(new_n508), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n515), .B2(G101), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT10), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n297), .B2(new_n299), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n521), .A2(new_n274), .B1(new_n509), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n513), .A2(new_n514), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT84), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n511), .A2(new_n512), .B1(new_n300), .B2(new_n509), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n287), .A3(new_n285), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n514), .A2(KEYINPUT12), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n531), .A2(KEYINPUT12), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G110), .B(G140), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n188), .A2(G227), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT79), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n514), .B1(new_n513), .B2(new_n524), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n527), .B2(new_n528), .ZN(new_n540));
  INV_X1    g354(.A(new_n537), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n534), .A2(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n488), .B1(new_n542), .B2(G469), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n529), .A2(new_n541), .A3(new_n533), .ZN(new_n544));
  INV_X1    g358(.A(new_n539), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n541), .B1(new_n529), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n487), .B(new_n242), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n486), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n300), .A2(new_n199), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n273), .B2(new_n199), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(G224), .A3(new_n188), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n188), .A2(G224), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n549), .B(new_n552), .C1(new_n273), .C2(new_n199), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT5), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n306), .B1(new_n311), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n555), .A2(new_n557), .B1(new_n315), .B2(new_n314), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n509), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n519), .A2(new_n520), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n317), .A2(new_n517), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT86), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n519), .A2(new_n520), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n317), .A2(new_n517), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n566), .A2(new_n567), .B1(new_n509), .B2(new_n558), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT86), .B1(new_n568), .B2(new_n560), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT6), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT85), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n560), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(KEYINPUT85), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(KEYINPUT6), .A3(new_n574), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n554), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n552), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n551), .A2(new_n553), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n563), .A2(new_n564), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n568), .A2(KEYINPUT86), .A3(new_n560), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n509), .A2(new_n558), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n509), .A2(new_n558), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n560), .B(KEYINPUT8), .Z(new_n588));
  OR2_X1    g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n550), .A2(new_n580), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n581), .A2(new_n584), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n242), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n578), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n582), .B2(new_n583), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n562), .B1(new_n519), .B2(new_n520), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n572), .B1(new_n598), .B2(new_n585), .ZN(new_n599));
  INV_X1    g413(.A(new_n560), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n599), .A2(new_n574), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n577), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n554), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n587), .A2(new_n588), .B1(new_n550), .B2(new_n580), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n582), .B2(new_n583), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n606), .B2(new_n581), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n593), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n595), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G214), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n385), .A2(new_n484), .A3(new_n548), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n604), .A2(new_n607), .A3(new_n615), .A4(new_n593), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n616), .A2(new_n610), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n594), .B1(new_n578), .B2(new_n592), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n604), .A2(new_n607), .A3(new_n593), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(KEYINPUT93), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n443), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n463), .A2(new_n472), .ZN(new_n624));
  INV_X1    g438(.A(new_n474), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n475), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(G478), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G478), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n242), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n626), .B2(new_n475), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n434), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n621), .A2(new_n622), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n342), .A2(new_n361), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n242), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n362), .B1(new_n643), .B2(G472), .ZN(new_n644));
  INV_X1    g458(.A(new_n254), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n548), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  AND2_X1   g463(.A1(new_n425), .A2(new_n427), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n650), .A2(new_n430), .B1(new_n428), .B2(KEYINPUT20), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n443), .B(KEYINPUT95), .Z(new_n652));
  NOR4_X1   g466(.A1(new_n651), .A2(new_n412), .A3(new_n482), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n617), .A2(new_n620), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n617), .A2(new_n620), .A3(new_n653), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT96), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n646), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT35), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  AND2_X1   g474(.A1(new_n252), .A2(new_n243), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n248), .A2(KEYINPUT77), .A3(new_n249), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n238), .B(new_n663), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n661), .A2(new_n662), .B1(new_n244), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n483), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n548), .A2(new_n666), .A3(new_n644), .A4(new_n612), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  INV_X1    g483(.A(new_n488), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n540), .A2(new_n541), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n529), .A2(new_n533), .ZN(new_n672));
  INV_X1    g486(.A(new_n538), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n671), .B(G469), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n547), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n486), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n664), .A2(new_n244), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n250), .B2(new_n253), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n256), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n363), .B1(new_n642), .B2(new_n680), .ZN(new_n681));
  AOI211_X1 g495(.A(KEYINPUT32), .B(new_n256), .C1(new_n342), .C2(new_n361), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n384), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n438), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n442), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n651), .A2(new_n412), .A3(new_n482), .A4(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n617), .A2(new_n620), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  INV_X1    g507(.A(KEYINPUT38), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n595), .B2(new_n608), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n595), .A2(new_n608), .A3(new_n694), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n370), .A2(new_n337), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n242), .B1(new_n379), .B2(new_n335), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n681), .B2(new_n682), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n434), .A2(new_n482), .A3(new_n611), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n698), .A2(new_n702), .A3(new_n665), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n688), .B(KEYINPUT39), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n548), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n258), .ZN(G45));
  NOR3_X1   g524(.A1(new_n434), .A2(new_n637), .A3(new_n689), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n617), .A2(new_n620), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n685), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  NAND3_X1  g528(.A1(new_n529), .A2(new_n541), .A3(new_n533), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n540), .B2(new_n541), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n242), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G469), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n718), .A2(new_n485), .A3(new_n547), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n385), .A2(new_n640), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND2_X1  g536(.A1(new_n657), .A2(new_n655), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n385), .A3(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  INV_X1    g539(.A(new_n621), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n683), .A2(new_n719), .A3(new_n726), .A4(new_n666), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  INV_X1    g542(.A(new_n652), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n485), .A3(new_n547), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n434), .A2(new_n482), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n617), .A2(new_n620), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n380), .A2(new_n335), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n256), .B1(new_n734), .B2(new_n361), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n643), .B2(G472), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT97), .B1(new_n736), .B2(new_n645), .ZN(new_n737));
  INV_X1    g551(.A(G472), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n642), .B2(new_n242), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT97), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n739), .A2(new_n254), .A3(new_n740), .A4(new_n735), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n733), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NOR3_X1   g557(.A1(new_n739), .A2(new_n665), .A3(new_n735), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n719), .A3(new_n726), .A4(new_n711), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  AOI21_X1  g560(.A(new_n738), .B1(new_n376), .B2(new_n382), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT100), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n367), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n681), .A2(new_n682), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT100), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n254), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n618), .A2(new_n485), .A3(new_n619), .A4(new_n610), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n529), .A2(new_n545), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n537), .ZN(new_n755));
  AOI21_X1  g569(.A(G902), .B1(new_n755), .B2(new_n715), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n488), .B1(new_n756), .B2(new_n487), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT98), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n672), .B2(new_n673), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n534), .A2(KEYINPUT98), .A3(new_n538), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n671), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n753), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n711), .A2(KEYINPUT42), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n752), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n683), .A2(new_n762), .A3(new_n645), .A4(new_n711), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n765), .A2(KEYINPUT99), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT99), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND3_X1  g584(.A1(new_n385), .A2(new_n690), .A3(new_n762), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  OAI21_X1  g586(.A(new_n678), .B1(new_n739), .B2(new_n362), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT102), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n632), .A2(new_n636), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n434), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT43), .Z(new_n777));
  AOI21_X1  g591(.A(KEYINPUT44), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n595), .A2(new_n608), .A3(new_n611), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n705), .A2(new_n485), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n487), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n671), .A4(new_n760), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n488), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n547), .B1(new_n787), .B2(KEYINPUT46), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n789), .B(new_n488), .C1(new_n785), .C2(new_n786), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n782), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT101), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT101), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(new_n782), .C1(new_n788), .C2(new_n790), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n773), .A2(KEYINPUT102), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n773), .A2(KEYINPUT102), .ZN(new_n797));
  OAI211_X1 g611(.A(KEYINPUT44), .B(new_n777), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(KEYINPUT103), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(KEYINPUT103), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n781), .B(new_n795), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  OAI21_X1  g616(.A(new_n485), .B1(new_n788), .B2(new_n790), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n485), .B(new_n804), .C1(new_n788), .C2(new_n790), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n779), .A2(new_n254), .A3(new_n711), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n683), .A2(KEYINPUT105), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT105), .B1(new_n683), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n806), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n200), .ZN(G42));
  XOR2_X1   g627(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n718), .A2(new_n547), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n442), .A3(new_n753), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n744), .A3(new_n777), .ZN(new_n818));
  INV_X1    g632(.A(new_n702), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n819), .A3(new_n645), .ZN(new_n820));
  INV_X1    g634(.A(new_n434), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n775), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n818), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n777), .A2(new_n441), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n736), .A2(new_n645), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n740), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n736), .A2(KEYINPUT97), .A3(new_n645), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n485), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n698), .A2(new_n831), .A3(new_n816), .A4(new_n610), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT50), .B1(new_n830), .B2(new_n832), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n825), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n816), .B(KEYINPUT107), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n486), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n785), .A2(new_n786), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n789), .B1(new_n838), .B2(new_n488), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n547), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n804), .B1(new_n841), .B2(new_n485), .ZN(new_n842));
  INV_X1    g656(.A(new_n807), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n830), .A2(new_n779), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n835), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(KEYINPUT112), .A3(new_n846), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n815), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n752), .A2(new_n777), .A3(new_n817), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT48), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n820), .A2(new_n639), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n440), .A3(G953), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n830), .A2(new_n726), .A3(new_n719), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n852), .A2(KEYINPUT48), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n830), .A2(new_n832), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n830), .A2(KEYINPUT50), .A3(new_n832), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n824), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n806), .A2(new_n807), .B1(new_n486), .B2(new_n836), .ZN(new_n865));
  OAI22_X1  g679(.A1(new_n864), .A2(KEYINPUT113), .B1(new_n865), .B2(new_n845), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT51), .B1(new_n835), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n859), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT114), .B1(new_n851), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n835), .A2(new_n867), .B1(new_n844), .B2(new_n846), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(KEYINPUT51), .C1(new_n867), .C2(new_n835), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n848), .B1(new_n865), .B2(new_n845), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n850), .A3(new_n864), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n814), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n859), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n610), .B(new_n729), .C1(new_n595), .C2(new_n608), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n412), .B(new_n482), .C1(new_n429), .C2(new_n433), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n638), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n645), .A3(new_n548), .A4(new_n644), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n645), .B1(new_n750), .B2(new_n747), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n548), .A2(new_n612), .A3(new_n484), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n882), .B(new_n667), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT108), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT108), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n613), .A2(new_n887), .A3(new_n667), .A4(new_n882), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n724), .A2(new_n742), .A3(new_n720), .A4(new_n727), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n482), .A2(new_n688), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n651), .A2(new_n892), .A3(new_n412), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n679), .A2(new_n683), .A3(new_n779), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n762), .A2(new_n744), .A3(new_n711), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n771), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n769), .A2(new_n889), .A3(new_n891), .A4(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n679), .B(new_n683), .C1(new_n691), .C2(new_n712), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n689), .A2(new_n831), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n620), .A2(new_n617), .A3(new_n731), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n757), .A2(new_n761), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n702), .A3(new_n665), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n745), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT109), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n904), .B(new_n906), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n890), .B1(new_n888), .B2(new_n886), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n769), .A4(new_n897), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n914));
  OAI22_X1  g728(.A1(new_n910), .A2(KEYINPUT53), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n910), .A2(KEYINPUT53), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n870), .A2(new_n877), .A3(new_n916), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n440), .A2(new_n188), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT115), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n836), .B(KEYINPUT49), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n696), .A2(new_n697), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n254), .A2(new_n486), .A3(new_n611), .A4(new_n776), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(KEYINPUT106), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(KEYINPUT106), .B2(new_n926), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n924), .A2(new_n819), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n929), .ZN(G75));
  NOR2_X1   g744(.A1(new_n188), .A2(G952), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n904), .B(KEYINPUT52), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n914), .B1(new_n898), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n765), .A2(new_n766), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT99), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n765), .A2(KEYINPUT99), .A3(new_n766), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n896), .B1(new_n939), .B2(new_n764), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n904), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT52), .B1(new_n904), .B2(KEYINPUT109), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n940), .A2(new_n943), .A3(KEYINPUT53), .A4(new_n912), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n242), .B1(new_n934), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT56), .B1(new_n945), .B2(G210), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n602), .B(KEYINPUT116), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n554), .B(KEYINPUT55), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n932), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n946), .B2(new_n950), .ZN(G51));
  NAND2_X1  g766(.A1(new_n934), .A2(new_n944), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n918), .B1(new_n934), .B2(new_n944), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n488), .B(KEYINPUT57), .Z(new_n957));
  OAI21_X1  g771(.A(new_n716), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n945), .A2(new_n838), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n931), .B1(new_n958), .B2(new_n959), .ZN(G54));
  AND3_X1   g774(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(new_n650), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n932), .B1(new_n961), .B2(new_n650), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G60));
  AND2_X1   g778(.A1(new_n630), .A2(new_n631), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n634), .B(KEYINPUT59), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n932), .B1(new_n956), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n919), .A2(new_n916), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n970), .B2(new_n967), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT117), .Z(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT60), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n934), .B2(new_n944), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n932), .B1(new_n977), .B2(new_n240), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n953), .A2(new_n664), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT118), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT118), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n977), .A2(new_n981), .A3(new_n664), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n978), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n977), .A2(new_n981), .A3(new_n664), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n981), .B1(new_n977), .B2(new_n664), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT119), .ZN(new_n987));
  INV_X1    g801(.A(new_n240), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n987), .B(new_n988), .C1(new_n917), .C2(new_n976), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT119), .B1(new_n977), .B2(new_n240), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI22_X1  g806(.A1(new_n983), .A2(KEYINPUT61), .B1(new_n986), .B2(new_n992), .ZN(G66));
  AOI21_X1  g807(.A(new_n188), .B1(new_n436), .B2(G224), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n912), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n947), .B1(G898), .B2(new_n188), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT120), .Z(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  INV_X1    g813(.A(KEYINPUT123), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n752), .A2(new_n726), .A3(new_n731), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n792), .B2(new_n794), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n812), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n899), .A2(new_n745), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n771), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n939), .B2(new_n764), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1003), .A2(new_n801), .A3(new_n188), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n369), .A2(new_n345), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT121), .Z(new_n1010));
  NAND2_X1  g824(.A1(new_n414), .A2(new_n416), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G900), .A2(G953), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT62), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1016), .B1(new_n709), .B2(new_n1004), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1005), .B(KEYINPUT62), .C1(new_n1020), .C2(new_n704), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n812), .ZN(new_n1023));
  INV_X1    g837(.A(new_n880), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n779), .B1(new_n1024), .B2(KEYINPUT122), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(KEYINPUT122), .B2(new_n1024), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n385), .A3(new_n706), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n801), .A2(new_n1022), .A3(new_n1023), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1028), .A2(G953), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1000), .B(new_n1015), .C1(new_n1029), .C2(new_n1012), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1015), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n801), .A2(new_n1022), .A3(new_n1023), .A4(new_n1027), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1012), .B1(new_n1032), .B2(new_n188), .ZN(new_n1033));
  OAI21_X1  g847(.A(KEYINPUT123), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1030), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1035), .ZN(new_n1037));
  OAI211_X1 g851(.A(KEYINPUT123), .B(new_n1037), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n1036), .A2(new_n1038), .ZN(G72));
  NAND2_X1  g853(.A1(new_n371), .A2(new_n374), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT126), .ZN(new_n1041));
  AOI22_X1  g855(.A1(new_n1040), .A2(new_n1041), .B1(new_n358), .B2(new_n359), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  NAND2_X1  g859(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT127), .Z(new_n1047));
  NAND2_X1  g861(.A1(new_n915), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1045), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1049), .B1(new_n1028), .B2(new_n912), .ZN(new_n1050));
  INV_X1    g864(.A(new_n699), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1003), .A2(new_n801), .A3(new_n912), .A4(new_n1007), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1053), .A2(KEYINPUT124), .A3(new_n1045), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n372), .A2(new_n335), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g870(.A(KEYINPUT124), .B1(new_n1053), .B2(new_n1045), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n932), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1058), .A2(KEYINPUT125), .ZN(new_n1059));
  INV_X1    g873(.A(KEYINPUT125), .ZN(new_n1060));
  OAI211_X1 g874(.A(new_n1060), .B(new_n932), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1052), .B1(new_n1059), .B2(new_n1061), .ZN(G57));
endmodule


