

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n796), .ZN(n780) );
  AND2_X1 U553 ( .A1(n779), .A2(n958), .ZN(n514) );
  NOR2_X1 U554 ( .A1(n733), .A2(n968), .ZN(n734) );
  AND2_X1 U555 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U556 ( .A(n725), .B(KEYINPUT96), .ZN(n728) );
  NAND2_X1 U557 ( .A1(n715), .A2(n714), .ZN(n750) );
  NOR2_X1 U558 ( .A1(G651), .A2(n635), .ZN(n655) );
  NOR2_X1 U559 ( .A1(n538), .A2(n537), .ZN(G160) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U561 ( .A1(n649), .A2(G89), .ZN(n515) );
  XNOR2_X1 U562 ( .A(n515), .B(KEYINPUT4), .ZN(n518) );
  XNOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .ZN(n516) );
  XNOR2_X1 U564 ( .A(n516), .B(KEYINPUT67), .ZN(n635) );
  INV_X1 U565 ( .A(G651), .ZN(n520) );
  NOR2_X1 U566 ( .A1(n635), .A2(n520), .ZN(n650) );
  NAND2_X1 U567 ( .A1(G76), .A2(n650), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U569 ( .A(n519), .B(KEYINPUT5), .ZN(n526) );
  NOR2_X1 U570 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n521), .Z(n654) );
  NAND2_X1 U572 ( .A1(G63), .A2(n654), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G51), .A2(n655), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U575 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n527), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U578 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n868) );
  NAND2_X1 U580 ( .A1(G113), .A2(n868), .ZN(n531) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XOR2_X1 U582 ( .A(KEYINPUT17), .B(n528), .Z(n529) );
  XNOR2_X2 U583 ( .A(KEYINPUT66), .B(n529), .ZN(n865) );
  NAND2_X1 U584 ( .A1(G137), .A2(n865), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n538) );
  INV_X1 U586 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n534), .A2(G2104), .ZN(n532) );
  XNOR2_X2 U588 ( .A(n532), .B(KEYINPUT65), .ZN(n864) );
  NAND2_X1 U589 ( .A1(G101), .A2(n864), .ZN(n533) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(n533), .Z(n536) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n534), .ZN(n870) );
  NAND2_X1 U592 ( .A1(n870), .A2(G125), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U594 ( .A1(G114), .A2(n868), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G126), .A2(n870), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G102), .A2(n864), .ZN(n541) );
  XOR2_X1 U598 ( .A(KEYINPUT85), .B(n541), .Z(n543) );
  NAND2_X1 U599 ( .A1(G138), .A2(n865), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U601 ( .A1(n545), .A2(n544), .ZN(G164) );
  XOR2_X1 U602 ( .A(G2443), .B(KEYINPUT102), .Z(n547) );
  XNOR2_X1 U603 ( .A(G2451), .B(G2427), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U605 ( .A(n548), .B(G2430), .Z(n550) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n549) );
  XNOR2_X1 U607 ( .A(n550), .B(n549), .ZN(n554) );
  XOR2_X1 U608 ( .A(KEYINPUT103), .B(G2438), .Z(n552) );
  XNOR2_X1 U609 ( .A(G2435), .B(G2454), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U611 ( .A(n554), .B(n553), .Z(n556) );
  XNOR2_X1 U612 ( .A(G2446), .B(KEYINPUT101), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n556), .B(n555), .ZN(n557) );
  AND2_X1 U614 ( .A1(n557), .A2(G14), .ZN(G401) );
  NAND2_X1 U615 ( .A1(G64), .A2(n654), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G52), .A2(n655), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G90), .A2(n649), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G77), .A2(n650), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U622 ( .A1(n564), .A2(n563), .ZN(G171) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  INV_X1 U626 ( .A(G82), .ZN(G220) );
  NAND2_X1 U627 ( .A1(n654), .A2(G62), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT83), .B(n565), .Z(n567) );
  NAND2_X1 U629 ( .A1(n655), .A2(G50), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT84), .B(n568), .Z(n572) );
  NAND2_X1 U632 ( .A1(G88), .A2(n649), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G75), .A2(n650), .ZN(n569) );
  AND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n819) );
  NAND2_X1 U639 ( .A1(n819), .A2(G567), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  XOR2_X1 U641 ( .A(G860), .B(KEYINPUT72), .Z(n607) );
  NAND2_X1 U642 ( .A1(G56), .A2(n654), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n575), .Z(n581) );
  NAND2_X1 U644 ( .A1(n649), .A2(G81), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G68), .A2(n650), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n655), .A2(G43), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n968) );
  OR2_X1 U652 ( .A1(n607), .A2(n968), .ZN(G153) );
  XNOR2_X1 U653 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n584), .B(KEYINPUT74), .ZN(n595) );
  INV_X1 U656 ( .A(G868), .ZN(n668) );
  NAND2_X1 U657 ( .A1(G54), .A2(n655), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT76), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G79), .A2(n650), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G66), .A2(n654), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G92), .A2(n649), .ZN(n588) );
  XNOR2_X1 U663 ( .A(KEYINPUT75), .B(n588), .ZN(n589) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n593), .Z(n969) );
  NAND2_X1 U667 ( .A1(n668), .A2(n969), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G78), .A2(n650), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n596), .B(KEYINPUT70), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G91), .A2(n649), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT69), .B(n597), .Z(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G65), .A2(n654), .ZN(n600) );
  XNOR2_X1 U675 ( .A(KEYINPUT71), .B(n600), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n655), .A2(G53), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G286), .A2(n668), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n607), .A2(G559), .ZN(n608) );
  INV_X1 U683 ( .A(n969), .ZN(n893) );
  NAND2_X1 U684 ( .A1(n608), .A2(n893), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U686 ( .A1(G559), .A2(n668), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n893), .A2(n610), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT77), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n968), .A2(G868), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G99), .A2(n864), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT78), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G111), .A2(n868), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G135), .A2(n865), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n870), .A2(G123), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT18), .B(n617), .Z(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U700 ( .A(KEYINPUT79), .B(n622), .ZN(n907) );
  XNOR2_X1 U701 ( .A(n907), .B(G2096), .ZN(n624) );
  INV_X1 U702 ( .A(G2100), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G93), .A2(n649), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G80), .A2(n650), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n655), .A2(G55), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT80), .B(n627), .Z(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n654), .A2(G67), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n667) );
  NAND2_X1 U712 ( .A1(G559), .A2(n893), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n968), .B(n632), .ZN(n665) );
  NOR2_X1 U714 ( .A1(n665), .A2(G860), .ZN(n633) );
  XNOR2_X1 U715 ( .A(n633), .B(KEYINPUT81), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n667), .B(n634), .ZN(G145) );
  NAND2_X1 U717 ( .A1(G87), .A2(n635), .ZN(n636) );
  XNOR2_X1 U718 ( .A(n636), .B(KEYINPUT82), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G49), .A2(n655), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U722 ( .A1(n654), .A2(n639), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(G288) );
  INV_X1 U724 ( .A(G303), .ZN(G166) );
  NAND2_X1 U725 ( .A1(G86), .A2(n649), .ZN(n643) );
  NAND2_X1 U726 ( .A1(G61), .A2(n654), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n650), .A2(G73), .ZN(n644) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U730 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n655), .A2(G48), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G85), .A2(n649), .ZN(n652) );
  NAND2_X1 U734 ( .A1(G72), .A2(n650), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U736 ( .A(KEYINPUT68), .B(n653), .Z(n659) );
  NAND2_X1 U737 ( .A1(G60), .A2(n654), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G47), .A2(n655), .ZN(n656) );
  AND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(G290) );
  XNOR2_X1 U741 ( .A(G288), .B(KEYINPUT19), .ZN(n661) );
  INV_X1 U742 ( .A(G299), .ZN(n956) );
  XNOR2_X1 U743 ( .A(n956), .B(G166), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n662), .B(G305), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n663), .B(n667), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n664), .B(G290), .ZN(n890) );
  XOR2_X1 U748 ( .A(n665), .B(n890), .Z(n666) );
  NAND2_X1 U749 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U760 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G96), .A2(n677), .ZN(n823) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n823), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G120), .A2(G108), .ZN(n678) );
  NOR2_X1 U764 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G69), .A2(n679), .ZN(n824) );
  NAND2_X1 U766 ( .A1(G567), .A2(n824), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n844) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U769 ( .A1(n844), .A2(n682), .ZN(n822) );
  NAND2_X1 U770 ( .A1(n822), .A2(G36), .ZN(G176) );
  XNOR2_X1 U771 ( .A(G1986), .B(KEYINPUT86), .ZN(n683) );
  XNOR2_X1 U772 ( .A(n683), .B(G290), .ZN(n966) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n715) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n715), .A2(n713), .ZN(n814) );
  NAND2_X1 U776 ( .A1(n966), .A2(n814), .ZN(n804) );
  NAND2_X1 U777 ( .A1(n864), .A2(G104), .ZN(n685) );
  NAND2_X1 U778 ( .A1(G140), .A2(n865), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U780 ( .A(KEYINPUT34), .B(n686), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G116), .A2(n868), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G128), .A2(n870), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U784 ( .A(KEYINPUT35), .B(n689), .Z(n690) );
  NOR2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U786 ( .A(KEYINPUT36), .B(n692), .ZN(n887) );
  XNOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NOR2_X1 U788 ( .A1(n887), .A2(n812), .ZN(n904) );
  NAND2_X1 U789 ( .A1(n814), .A2(n904), .ZN(n810) );
  NAND2_X1 U790 ( .A1(G119), .A2(n870), .ZN(n694) );
  NAND2_X1 U791 ( .A1(G131), .A2(n865), .ZN(n693) );
  NAND2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G107), .A2(n868), .ZN(n696) );
  NAND2_X1 U794 ( .A1(G95), .A2(n864), .ZN(n695) );
  NAND2_X1 U795 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U796 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U797 ( .A(n699), .B(KEYINPUT87), .ZN(n859) );
  AND2_X1 U798 ( .A1(n859), .A2(G1991), .ZN(n710) );
  XOR2_X1 U799 ( .A(KEYINPUT89), .B(KEYINPUT38), .Z(n701) );
  NAND2_X1 U800 ( .A1(G105), .A2(n864), .ZN(n700) );
  XNOR2_X1 U801 ( .A(n701), .B(n700), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G129), .A2(n870), .ZN(n703) );
  NAND2_X1 U803 ( .A1(G141), .A2(n865), .ZN(n702) );
  NAND2_X1 U804 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U805 ( .A1(n868), .A2(G117), .ZN(n704) );
  XOR2_X1 U806 ( .A(KEYINPUT88), .B(n704), .Z(n705) );
  NOR2_X1 U807 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n881) );
  AND2_X1 U809 ( .A1(n881), .A2(G1996), .ZN(n709) );
  NOR2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n909) );
  INV_X1 U811 ( .A(n814), .ZN(n711) );
  NOR2_X1 U812 ( .A1(n909), .A2(n711), .ZN(n807) );
  INV_X1 U813 ( .A(n807), .ZN(n712) );
  NAND2_X1 U814 ( .A1(n810), .A2(n712), .ZN(n802) );
  INV_X1 U815 ( .A(n713), .ZN(n714) );
  BUF_X1 U816 ( .A(n750), .Z(n761) );
  XNOR2_X1 U817 ( .A(G1961), .B(KEYINPUT91), .ZN(n1002) );
  NAND2_X1 U818 ( .A1(n761), .A2(n1002), .ZN(n716) );
  XNOR2_X1 U819 ( .A(n716), .B(KEYINPUT92), .ZN(n719) );
  INV_X1 U820 ( .A(n750), .ZN(n735) );
  XOR2_X1 U821 ( .A(G2078), .B(KEYINPUT25), .Z(n717) );
  XNOR2_X1 U822 ( .A(KEYINPUT93), .B(n717), .ZN(n930) );
  NAND2_X1 U823 ( .A1(n735), .A2(n930), .ZN(n718) );
  NAND2_X1 U824 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U825 ( .A(KEYINPUT94), .B(n720), .ZN(n755) );
  NAND2_X1 U826 ( .A1(G171), .A2(n755), .ZN(n721) );
  XOR2_X1 U827 ( .A(KEYINPUT95), .B(n721), .Z(n749) );
  NAND2_X1 U828 ( .A1(n735), .A2(G2072), .ZN(n722) );
  XOR2_X1 U829 ( .A(KEYINPUT27), .B(n722), .Z(n724) );
  NAND2_X1 U830 ( .A1(G1956), .A2(n761), .ZN(n723) );
  NOR2_X1 U831 ( .A1(n956), .A2(n728), .ZN(n727) );
  XNOR2_X1 U832 ( .A(KEYINPUT28), .B(KEYINPUT97), .ZN(n726) );
  XNOR2_X1 U833 ( .A(n727), .B(n726), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n956), .A2(n728), .ZN(n744) );
  INV_X1 U835 ( .A(G1996), .ZN(n931) );
  NOR2_X1 U836 ( .A1(n750), .A2(n931), .ZN(n730) );
  XOR2_X1 U837 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n729) );
  XNOR2_X1 U838 ( .A(n730), .B(n729), .ZN(n732) );
  NAND2_X1 U839 ( .A1(n750), .A2(G1341), .ZN(n731) );
  NAND2_X1 U840 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U841 ( .A(n734), .B(KEYINPUT64), .Z(n740) );
  OR2_X1 U842 ( .A1(n740), .A2(n969), .ZN(n739) );
  NOR2_X1 U843 ( .A1(n735), .A2(G1348), .ZN(n737) );
  NOR2_X1 U844 ( .A1(G2067), .A2(n761), .ZN(n736) );
  NOR2_X1 U845 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U846 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U847 ( .A1(n740), .A2(n969), .ZN(n741) );
  NAND2_X1 U848 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U849 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U850 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U851 ( .A(KEYINPUT29), .B(n747), .Z(n748) );
  NAND2_X1 U852 ( .A1(n749), .A2(n748), .ZN(n760) );
  NAND2_X1 U853 ( .A1(G8), .A2(n750), .ZN(n796) );
  NOR2_X1 U854 ( .A1(G1966), .A2(n796), .ZN(n772) );
  NOR2_X1 U855 ( .A1(G2084), .A2(n761), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n772), .A2(n769), .ZN(n751) );
  XOR2_X1 U857 ( .A(KEYINPUT99), .B(n751), .Z(n752) );
  NAND2_X1 U858 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U859 ( .A(KEYINPUT30), .B(n753), .ZN(n754) );
  NOR2_X1 U860 ( .A1(G168), .A2(n754), .ZN(n757) );
  NOR2_X1 U861 ( .A1(G171), .A2(n755), .ZN(n756) );
  NOR2_X1 U862 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U863 ( .A(KEYINPUT31), .B(n758), .Z(n759) );
  NAND2_X1 U864 ( .A1(n760), .A2(n759), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n770), .A2(G286), .ZN(n766) );
  NOR2_X1 U866 ( .A1(G1971), .A2(n796), .ZN(n763) );
  NOR2_X1 U867 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U868 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U869 ( .A1(n764), .A2(G303), .ZN(n765) );
  NAND2_X1 U870 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U871 ( .A1(G8), .A2(n767), .ZN(n768) );
  XNOR2_X1 U872 ( .A(n768), .B(KEYINPUT32), .ZN(n776) );
  NAND2_X1 U873 ( .A1(G8), .A2(n769), .ZN(n774) );
  INV_X1 U874 ( .A(n770), .ZN(n771) );
  NOR2_X1 U875 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U876 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U877 ( .A1(n776), .A2(n775), .ZN(n790) );
  NOR2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n957) );
  NOR2_X1 U879 ( .A1(G1971), .A2(G303), .ZN(n777) );
  NOR2_X1 U880 ( .A1(n957), .A2(n777), .ZN(n778) );
  NAND2_X1 U881 ( .A1(n790), .A2(n778), .ZN(n779) );
  NAND2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NAND2_X1 U883 ( .A1(n514), .A2(n780), .ZN(n782) );
  INV_X1 U884 ( .A(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U885 ( .A1(n782), .A2(n781), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n957), .A2(KEYINPUT33), .ZN(n783) );
  NOR2_X1 U887 ( .A1(n783), .A2(n796), .ZN(n785) );
  XOR2_X1 U888 ( .A(G1981), .B(G305), .Z(n953) );
  INV_X1 U889 ( .A(n953), .ZN(n784) );
  NOR2_X1 U890 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U891 ( .A1(n787), .A2(n786), .ZN(n800) );
  NOR2_X1 U892 ( .A1(G2090), .A2(G303), .ZN(n788) );
  XNOR2_X1 U893 ( .A(n788), .B(KEYINPUT100), .ZN(n789) );
  NAND2_X1 U894 ( .A1(n789), .A2(G8), .ZN(n791) );
  NAND2_X1 U895 ( .A1(n791), .A2(n790), .ZN(n792) );
  AND2_X1 U896 ( .A1(n792), .A2(n796), .ZN(n798) );
  NOR2_X1 U897 ( .A1(G1981), .A2(G305), .ZN(n793) );
  XOR2_X1 U898 ( .A(n793), .B(KEYINPUT24), .Z(n794) );
  XNOR2_X1 U899 ( .A(KEYINPUT90), .B(n794), .ZN(n795) );
  NOR2_X1 U900 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U901 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U902 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U903 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U904 ( .A1(n804), .A2(n803), .ZN(n817) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n881), .ZN(n919) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n859), .ZN(n911) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U908 ( .A1(n911), .A2(n805), .ZN(n806) );
  NOR2_X1 U909 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U910 ( .A1(n919), .A2(n808), .ZN(n809) );
  XNOR2_X1 U911 ( .A(n809), .B(KEYINPUT39), .ZN(n811) );
  NAND2_X1 U912 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U913 ( .A1(n887), .A2(n812), .ZN(n903) );
  NAND2_X1 U914 ( .A1(n813), .A2(n903), .ZN(n815) );
  NAND2_X1 U915 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U920 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U922 ( .A1(n822), .A2(n821), .ZN(G188) );
  NOR2_X1 U923 ( .A1(n824), .A2(n823), .ZN(G325) );
  XOR2_X1 U924 ( .A(KEYINPUT104), .B(G325), .Z(G261) );
  XOR2_X1 U925 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  XOR2_X1 U929 ( .A(G2100), .B(G2096), .Z(n826) );
  XNOR2_X1 U930 ( .A(KEYINPUT42), .B(G2678), .ZN(n825) );
  XNOR2_X1 U931 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U932 ( .A(KEYINPUT43), .B(G2090), .Z(n828) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n827) );
  XNOR2_X1 U934 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U935 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n831) );
  XNOR2_X1 U937 ( .A(n832), .B(n831), .ZN(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT107), .B(G1976), .Z(n834) );
  XNOR2_X1 U939 ( .A(G1956), .B(G1961), .ZN(n833) );
  XNOR2_X1 U940 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U941 ( .A(n835), .B(KEYINPUT41), .Z(n837) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U943 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U944 ( .A(G1981), .B(G1971), .Z(n839) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U946 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U947 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U948 ( .A(KEYINPUT106), .B(G2474), .ZN(n842) );
  XNOR2_X1 U949 ( .A(n843), .B(n842), .ZN(G229) );
  XNOR2_X1 U950 ( .A(KEYINPUT105), .B(n844), .ZN(G319) );
  NAND2_X1 U951 ( .A1(n870), .A2(G124), .ZN(n845) );
  XNOR2_X1 U952 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U953 ( .A1(G100), .A2(n864), .ZN(n846) );
  NAND2_X1 U954 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U955 ( .A1(G112), .A2(n868), .ZN(n849) );
  NAND2_X1 U956 ( .A1(G136), .A2(n865), .ZN(n848) );
  NAND2_X1 U957 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U958 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G118), .A2(n868), .ZN(n853) );
  NAND2_X1 U960 ( .A1(G130), .A2(n870), .ZN(n852) );
  NAND2_X1 U961 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n864), .A2(G106), .ZN(n855) );
  NAND2_X1 U963 ( .A1(G142), .A2(n865), .ZN(n854) );
  NAND2_X1 U964 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U965 ( .A(n856), .B(KEYINPUT45), .Z(n857) );
  NOR2_X1 U966 ( .A1(n858), .A2(n857), .ZN(n860) );
  XNOR2_X1 U967 ( .A(n860), .B(n859), .ZN(n880) );
  XOR2_X1 U968 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n862) );
  XNOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n861) );
  XNOR2_X1 U970 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U971 ( .A(n863), .B(KEYINPUT113), .Z(n878) );
  NAND2_X1 U972 ( .A1(n864), .A2(G103), .ZN(n867) );
  NAND2_X1 U973 ( .A1(G139), .A2(n865), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n867), .A2(n866), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n868), .A2(G115), .ZN(n869) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(n869), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n870), .A2(G127), .ZN(n871) );
  XOR2_X1 U978 ( .A(KEYINPUT110), .B(n871), .Z(n872) );
  NOR2_X1 U979 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U980 ( .A(n874), .B(KEYINPUT47), .ZN(n875) );
  NOR2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n914) );
  XNOR2_X1 U982 ( .A(n914), .B(KEYINPUT48), .ZN(n877) );
  XNOR2_X1 U983 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U984 ( .A(n880), .B(n879), .Z(n883) );
  XOR2_X1 U985 ( .A(G164), .B(n881), .Z(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(n884), .B(n907), .Z(n886) );
  XNOR2_X1 U988 ( .A(G160), .B(G162), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U990 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U991 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n968), .B(G171), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U996 ( .A1(G37), .A2(n895), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n896) );
  XOR2_X1 U998 ( .A(KEYINPUT114), .B(n896), .Z(n897) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n897), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n898) );
  XOR2_X1 U1001 ( .A(KEYINPUT115), .B(n898), .Z(n899) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n899), .ZN(n900) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n900), .ZN(n901) );
  NAND2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  INV_X1 U1007 ( .A(n903), .ZN(n905) );
  NOR2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n913) );
  XOR2_X1 U1009 ( .A(G2084), .B(G160), .Z(n906) );
  NOR2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n924) );
  XOR2_X1 U1014 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT50), .B(n917), .ZN(n922) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n920), .Z(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT52), .B(n925), .ZN(n926) );
  INV_X1 U1024 ( .A(KEYINPUT55), .ZN(n949) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n949), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(G29), .ZN(n1013) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(G2090), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(G35), .ZN(n947) );
  XNOR2_X1 U1029 ( .A(G2084), .B(G34), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(KEYINPUT54), .ZN(n945) );
  XNOR2_X1 U1031 ( .A(G27), .B(n930), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(G32), .B(n931), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(n932), .A2(G28), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G25), .B(G1991), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT118), .B(n933), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(G2072), .B(G33), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(n940), .B(KEYINPUT119), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT53), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n949), .B(n948), .ZN(n951) );
  INV_X1 U1047 ( .A(G29), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n952), .ZN(n1011) );
  XNOR2_X1 U1050 ( .A(G16), .B(KEYINPUT56), .ZN(n982) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(KEYINPUT57), .B(n955), .ZN(n980) );
  XNOR2_X1 U1054 ( .A(n956), .B(G1956), .ZN(n964) );
  XOR2_X1 U1055 ( .A(n957), .B(KEYINPUT122), .Z(n959) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1057 ( .A(G1971), .B(G303), .Z(n960) );
  XNOR2_X1 U1058 ( .A(KEYINPUT123), .B(n960), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT124), .B(n967), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(n968), .B(G1341), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT120), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(n969), .ZN(n972) );
  XOR2_X1 U1066 ( .A(G171), .B(G1961), .Z(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT121), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(KEYINPUT125), .B(n978), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n1009) );
  INV_X1 U1074 ( .A(G16), .ZN(n1007) );
  XNOR2_X1 U1075 ( .A(KEYINPUT127), .B(G1966), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(G21), .ZN(n1001) );
  XNOR2_X1 U1077 ( .A(G1341), .B(G19), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G6), .B(G1981), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n991) );
  XOR2_X1 U1080 ( .A(KEYINPUT126), .B(G4), .Z(n987) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(n987), .B(n986), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G1956), .B(G20), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT60), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n994) );
  XNOR2_X1 U1088 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n996) );
  XOR2_X1 U1090 ( .A(G1986), .B(G24), .Z(n995) );
  NAND2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n997), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1095 ( .A(G5), .B(n1002), .Z(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(KEYINPUT61), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1014), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

