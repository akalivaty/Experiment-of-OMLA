

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744;

  OR2_X1 U378 ( .A1(n387), .A2(n648), .ZN(n382) );
  INV_X1 U379 ( .A(n645), .ZN(n387) );
  XNOR2_X1 U380 ( .A(n570), .B(KEYINPUT77), .ZN(n586) );
  AND2_X2 U381 ( .A1(n597), .A2(n598), .ZN(n390) );
  XNOR2_X2 U382 ( .A(G143), .B(G128), .ZN(n481) );
  XNOR2_X2 U383 ( .A(n594), .B(KEYINPUT19), .ZN(n576) );
  NAND2_X2 U384 ( .A1(n584), .A2(n681), .ZN(n594) );
  XNOR2_X2 U385 ( .A(n472), .B(KEYINPUT16), .ZN(n717) );
  NOR2_X1 U386 ( .A1(n540), .A2(n539), .ZN(n648) );
  NOR2_X1 U387 ( .A1(n523), .A2(n599), .ZN(n537) );
  NOR2_X1 U388 ( .A1(n739), .A2(n744), .ZN(n575) );
  XNOR2_X1 U389 ( .A(n382), .B(KEYINPUT99), .ZN(n686) );
  NOR2_X1 U390 ( .A1(n422), .A2(n426), .ZN(n631) );
  NOR2_X1 U391 ( .A1(n627), .A2(n711), .ZN(n383) );
  NOR2_X1 U392 ( .A1(n703), .A2(n711), .ZN(n389) );
  NOR2_X1 U393 ( .A1(n619), .A2(n711), .ZN(n621) );
  NOR2_X1 U394 ( .A1(n710), .A2(n711), .ZN(n393) );
  NAND2_X1 U395 ( .A1(n425), .A2(n423), .ZN(n422) );
  AND2_X1 U396 ( .A1(n537), .A2(n366), .ZN(n639) );
  AND2_X1 U397 ( .A1(n432), .A2(n431), .ZN(n577) );
  XNOR2_X1 U398 ( .A(n550), .B(n549), .ZN(n558) );
  NOR2_X1 U399 ( .A1(n685), .A2(n684), .ZN(n550) );
  NOR2_X1 U400 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U401 ( .A(n557), .B(n418), .ZN(n599) );
  XNOR2_X1 U402 ( .A(n505), .B(n504), .ZN(n540) );
  XNOR2_X1 U403 ( .A(n381), .B(n497), .ZN(n622) );
  XNOR2_X1 U404 ( .A(n439), .B(n399), .ZN(n454) );
  BUF_X1 U405 ( .A(n720), .Z(n355) );
  XNOR2_X1 U406 ( .A(n374), .B(G101), .ZN(n473) );
  XNOR2_X1 U407 ( .A(n437), .B(G116), .ZN(n471) );
  XNOR2_X1 U408 ( .A(G137), .B(G140), .ZN(n511) );
  INV_X2 U409 ( .A(KEYINPUT3), .ZN(n421) );
  NOR2_X1 U410 ( .A1(n707), .A2(n364), .ZN(n426) );
  XNOR2_X1 U411 ( .A(n444), .B(n445), .ZN(n726) );
  XNOR2_X1 U412 ( .A(n726), .B(n356), .ZN(n510) );
  XNOR2_X1 U413 ( .A(n435), .B(G146), .ZN(n476) );
  INV_X1 U414 ( .A(G125), .ZN(n435) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n495) );
  XNOR2_X1 U416 ( .A(n478), .B(n498), .ZN(n444) );
  XNOR2_X1 U417 ( .A(G902), .B(KEYINPUT15), .ZN(n483) );
  XNOR2_X1 U418 ( .A(n555), .B(KEYINPUT69), .ZN(n591) );
  XNOR2_X1 U419 ( .A(G469), .B(n517), .ZN(n557) );
  INV_X1 U420 ( .A(G472), .ZN(n386) );
  XNOR2_X1 U421 ( .A(G478), .B(KEYINPUT98), .ZN(n506) );
  NAND2_X1 U422 ( .A1(n643), .A2(n587), .ZN(n376) );
  XOR2_X1 U423 ( .A(KEYINPUT93), .B(G110), .Z(n459) );
  XNOR2_X1 U424 ( .A(G128), .B(G119), .ZN(n458) );
  XNOR2_X1 U425 ( .A(n398), .B(n396), .ZN(n457) );
  XNOR2_X1 U426 ( .A(n511), .B(n397), .ZN(n396) );
  NAND2_X1 U427 ( .A1(n454), .A2(G221), .ZN(n398) );
  XNOR2_X1 U428 ( .A(n455), .B(KEYINPUT85), .ZN(n397) );
  XNOR2_X1 U429 ( .A(G122), .B(G143), .ZN(n499) );
  XNOR2_X1 U430 ( .A(n476), .B(n434), .ZN(n728) );
  INV_X1 U431 ( .A(KEYINPUT10), .ZN(n434) );
  INV_X1 U432 ( .A(G107), .ZN(n513) );
  XNOR2_X1 U433 ( .A(n512), .B(n414), .ZN(n725) );
  INV_X1 U434 ( .A(KEYINPUT92), .ZN(n414) );
  XOR2_X1 U435 ( .A(n510), .B(n451), .Z(n630) );
  XNOR2_X1 U436 ( .A(G110), .B(G104), .ZN(n719) );
  XNOR2_X1 U437 ( .A(KEYINPUT17), .B(KEYINPUT79), .ZN(n394) );
  XNOR2_X1 U438 ( .A(n378), .B(n477), .ZN(n479) );
  XNOR2_X1 U439 ( .A(n473), .B(n373), .ZN(n474) );
  XNOR2_X1 U440 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U441 ( .A(KEYINPUT102), .ZN(n416) );
  INV_X1 U442 ( .A(KEYINPUT1), .ZN(n418) );
  XNOR2_X1 U443 ( .A(n571), .B(KEYINPUT39), .ZN(n572) );
  INV_X1 U444 ( .A(KEYINPUT87), .ZN(n571) );
  AND2_X1 U445 ( .A1(n388), .A2(n387), .ZN(n593) );
  XNOR2_X1 U446 ( .A(n592), .B(KEYINPUT103), .ZN(n388) );
  INV_X1 U447 ( .A(n599), .ZN(n666) );
  XNOR2_X1 U448 ( .A(n465), .B(n464), .ZN(n520) );
  XNOR2_X1 U449 ( .A(n463), .B(KEYINPUT25), .ZN(n464) );
  INV_X1 U450 ( .A(n453), .ZN(n675) );
  INV_X1 U451 ( .A(n520), .ZN(n669) );
  NAND2_X1 U452 ( .A1(n412), .A2(n411), .ZN(n410) );
  XNOR2_X1 U453 ( .A(n471), .B(n369), .ZN(n442) );
  XNOR2_X1 U454 ( .A(n438), .B(KEYINPUT7), .ZN(n369) );
  INV_X1 U455 ( .A(KEYINPUT83), .ZN(n375) );
  INV_X1 U456 ( .A(KEYINPUT24), .ZN(n455) );
  XOR2_X1 U457 ( .A(G104), .B(G113), .Z(n500) );
  XNOR2_X1 U458 ( .A(n371), .B(n370), .ZN(n596) );
  INV_X1 U459 ( .A(KEYINPUT72), .ZN(n370) );
  NOR2_X1 U460 ( .A1(n589), .A2(n588), .ZN(n371) );
  XNOR2_X1 U461 ( .A(n376), .B(n375), .ZN(n588) );
  NOR2_X1 U462 ( .A1(n357), .A2(KEYINPUT76), .ZN(n403) );
  INV_X1 U463 ( .A(KEYINPUT8), .ZN(n399) );
  INV_X1 U464 ( .A(KEYINPUT67), .ZN(n374) );
  INV_X1 U465 ( .A(KEYINPUT78), .ZN(n373) );
  XNOR2_X1 U466 ( .A(n478), .B(n358), .ZN(n378) );
  OR2_X1 U467 ( .A1(G902), .A2(G237), .ZN(n486) );
  NAND2_X1 U468 ( .A1(n539), .A2(n531), .ZN(n684) );
  XNOR2_X1 U469 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n461) );
  AND2_X1 U470 ( .A1(n599), .A2(n417), .ZN(n541) );
  INV_X1 U471 ( .A(n665), .ZN(n417) );
  NAND2_X1 U472 ( .A1(n520), .A2(n400), .ZN(n665) );
  XNOR2_X1 U473 ( .A(n379), .B(n456), .ZN(n616) );
  XNOR2_X1 U474 ( .A(n457), .B(n460), .ZN(n379) );
  XOR2_X1 U475 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n438) );
  XNOR2_X1 U476 ( .A(G107), .B(G122), .ZN(n437) );
  XNOR2_X1 U477 ( .A(n503), .B(n496), .ZN(n381) );
  XNOR2_X1 U478 ( .A(n413), .B(n510), .ZN(n704) );
  XNOR2_X1 U479 ( .A(n415), .B(n725), .ZN(n413) );
  INV_X1 U480 ( .A(n558), .ZN(n680) );
  XNOR2_X1 U481 ( .A(n433), .B(n556), .ZN(n432) );
  NOR2_X1 U482 ( .A1(n665), .A2(n557), .ZN(n561) );
  XNOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT0), .ZN(n489) );
  AND2_X1 U484 ( .A1(n552), .A2(n488), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n562), .B(n362), .ZN(n590) );
  NAND2_X1 U486 ( .A1(n707), .A2(n365), .ZN(n425) );
  NOR2_X1 U487 ( .A1(n424), .A2(n711), .ZN(n423) );
  NOR2_X1 U488 ( .A1(n364), .A2(G472), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n516), .B(n394), .ZN(n480) );
  XNOR2_X1 U490 ( .A(n395), .B(n363), .ZN(n739) );
  NOR2_X1 U491 ( .A1(n384), .A2(n666), .ZN(n651) );
  XNOR2_X1 U492 ( .A(n595), .B(n385), .ZN(n384) );
  INV_X1 U493 ( .A(KEYINPUT36), .ZN(n385) );
  INV_X1 U494 ( .A(KEYINPUT35), .ZN(n532) );
  NAND2_X1 U495 ( .A1(n540), .A2(n539), .ZN(n645) );
  NOR2_X1 U496 ( .A1(n675), .A2(n367), .ZN(n366) );
  XNOR2_X1 U497 ( .A(n612), .B(n391), .ZN(n614) );
  INV_X1 U498 ( .A(n613), .ZN(n391) );
  INV_X1 U499 ( .A(n668), .ZN(n400) );
  XOR2_X1 U500 ( .A(n473), .B(G146), .Z(n356) );
  AND2_X1 U501 ( .A1(n656), .A2(n654), .ZN(n357) );
  AND2_X1 U502 ( .A1(G224), .A2(n720), .ZN(n358) );
  AND2_X1 U503 ( .A1(n508), .A2(n400), .ZN(n359) );
  AND2_X1 U504 ( .A1(n357), .A2(KEYINPUT76), .ZN(n360) );
  XNOR2_X1 U505 ( .A(n509), .B(KEYINPUT22), .ZN(n361) );
  XOR2_X1 U506 ( .A(KEYINPUT6), .B(KEYINPUT100), .Z(n362) );
  XOR2_X1 U507 ( .A(n574), .B(KEYINPUT40), .Z(n363) );
  XOR2_X1 U508 ( .A(n630), .B(n629), .Z(n364) );
  AND2_X1 U509 ( .A1(n364), .A2(G472), .ZN(n365) );
  INV_X1 U510 ( .A(G953), .ZN(n720) );
  NOR2_X1 U511 ( .A1(G952), .A2(n355), .ZN(n711) );
  INV_X1 U512 ( .A(n711), .ZN(n427) );
  INV_X1 U513 ( .A(n669), .ZN(n367) );
  NOR2_X1 U514 ( .A1(n368), .A2(n644), .ZN(n580) );
  XNOR2_X1 U515 ( .A(n579), .B(n578), .ZN(n368) );
  XNOR2_X1 U516 ( .A(n573), .B(n572), .ZN(n606) );
  XNOR2_X1 U517 ( .A(n717), .B(n372), .ZN(n377) );
  XNOR2_X1 U518 ( .A(n475), .B(n479), .ZN(n372) );
  NOR2_X1 U519 ( .A1(n605), .A2(KEYINPUT76), .ZN(n404) );
  XNOR2_X1 U520 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U521 ( .A(n377), .B(n482), .ZN(n700) );
  NOR2_X1 U522 ( .A1(n639), .A2(n743), .ZN(n525) );
  NAND2_X1 U523 ( .A1(n591), .A2(n675), .ZN(n433) );
  NAND2_X1 U524 ( .A1(n707), .A2(G469), .ZN(n708) );
  XNOR2_X2 U525 ( .A(n380), .B(n361), .ZN(n523) );
  NAND2_X1 U526 ( .A1(n543), .A2(n359), .ZN(n380) );
  XNOR2_X1 U527 ( .A(n442), .B(n441), .ZN(n613) );
  XNOR2_X1 U528 ( .A(n541), .B(n416), .ZN(n527) );
  XNOR2_X1 U529 ( .A(n516), .B(n515), .ZN(n415) );
  NOR2_X1 U530 ( .A1(n690), .A2(n530), .ZN(n408) );
  XNOR2_X1 U531 ( .A(n529), .B(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U532 ( .A1(n404), .A2(n403), .ZN(n402) );
  XNOR2_X1 U533 ( .A(n383), .B(n628), .ZN(G60) );
  XNOR2_X2 U534 ( .A(n452), .B(n386), .ZN(n562) );
  XNOR2_X1 U535 ( .A(n389), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X2 U536 ( .A(n390), .B(KEYINPUT48), .ZN(n605) );
  NAND2_X1 U537 ( .A1(n402), .A2(n401), .ZN(n405) );
  NAND2_X1 U538 ( .A1(n392), .A2(n740), .ZN(n535) );
  XNOR2_X1 U539 ( .A(n525), .B(n526), .ZN(n392) );
  XNOR2_X1 U540 ( .A(n393), .B(KEYINPUT118), .ZN(G54) );
  NAND2_X1 U541 ( .A1(n576), .A2(n429), .ZN(n428) );
  NAND2_X1 U542 ( .A1(n606), .A2(n387), .ZN(n395) );
  AND2_X1 U543 ( .A1(n605), .A2(n357), .ZN(n730) );
  NAND2_X1 U544 ( .A1(n605), .A2(n360), .ZN(n401) );
  NAND2_X1 U545 ( .A1(n605), .A2(n656), .ZN(n611) );
  NAND2_X1 U546 ( .A1(n405), .A2(n712), .ZN(n412) );
  XNOR2_X2 U547 ( .A(n406), .B(n532), .ZN(n740) );
  NAND2_X1 U548 ( .A1(n407), .A2(n583), .ZN(n406) );
  XNOR2_X1 U549 ( .A(n408), .B(KEYINPUT34), .ZN(n407) );
  AND2_X4 U550 ( .A1(n409), .A2(n410), .ZN(n707) );
  AND2_X2 U551 ( .A1(n659), .A2(n610), .ZN(n409) );
  NAND2_X1 U552 ( .A1(n712), .A2(n609), .ZN(n659) );
  INV_X1 U553 ( .A(KEYINPUT2), .ZN(n411) );
  XOR2_X2 U554 ( .A(KEYINPUT68), .B(G131), .Z(n498) );
  XNOR2_X2 U555 ( .A(n420), .B(n419), .ZN(n470) );
  XNOR2_X2 U556 ( .A(G113), .B(G119), .ZN(n419) );
  XNOR2_X2 U557 ( .A(n421), .B(KEYINPUT90), .ZN(n420) );
  NOR2_X1 U558 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X2 U559 ( .A(n428), .B(n489), .ZN(n543) );
  XNOR2_X2 U560 ( .A(n430), .B(KEYINPUT45), .ZN(n712) );
  NAND2_X1 U561 ( .A1(n548), .A2(n547), .ZN(n430) );
  INV_X1 U562 ( .A(n557), .ZN(n431) );
  NAND2_X1 U563 ( .A1(n614), .A2(n427), .ZN(n615) );
  INV_X1 U564 ( .A(n540), .ZN(n531) );
  XOR2_X2 U565 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n478) );
  XNOR2_X1 U566 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n436) );
  INV_X1 U567 ( .A(KEYINPUT74), .ZN(n578) );
  XNOR2_X1 U568 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U569 ( .A(n474), .B(KEYINPUT18), .ZN(n475) );
  XNOR2_X1 U570 ( .A(n563), .B(KEYINPUT107), .ZN(n564) );
  XNOR2_X1 U571 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n445), .B(n440), .ZN(n441) );
  INV_X1 U573 ( .A(KEYINPUT109), .ZN(n574) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n539) );
  INV_X1 U575 ( .A(KEYINPUT123), .ZN(n620) );
  XNOR2_X1 U576 ( .A(n615), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U577 ( .A(G134), .B(n481), .ZN(n445) );
  NAND2_X1 U578 ( .A1(n720), .A2(G234), .ZN(n439) );
  NAND2_X1 U579 ( .A1(G217), .A2(n454), .ZN(n440) );
  INV_X1 U580 ( .A(n483), .ZN(n610) );
  INV_X1 U581 ( .A(KEYINPUT44), .ZN(n443) );
  NAND2_X1 U582 ( .A1(n443), .A2(KEYINPUT88), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n447) );
  XNOR2_X1 U584 ( .A(G116), .B(G137), .ZN(n446) );
  XNOR2_X1 U585 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U586 ( .A(n448), .B(n470), .Z(n450) );
  NAND2_X1 U587 ( .A1(n495), .A2(G210), .ZN(n449) );
  XNOR2_X1 U588 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U589 ( .A1(n630), .A2(G902), .ZN(n452) );
  INV_X1 U590 ( .A(n562), .ZN(n453) );
  XNOR2_X1 U591 ( .A(n728), .B(KEYINPUT23), .ZN(n456) );
  XNOR2_X1 U592 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U593 ( .A1(n616), .A2(G902), .ZN(n465) );
  NAND2_X1 U594 ( .A1(n483), .A2(G234), .ZN(n462) );
  XNOR2_X1 U595 ( .A(n462), .B(n461), .ZN(n490) );
  NAND2_X1 U596 ( .A1(G217), .A2(n490), .ZN(n463) );
  NAND2_X1 U597 ( .A1(G237), .A2(G234), .ZN(n466) );
  XNOR2_X1 U598 ( .A(n466), .B(KEYINPUT14), .ZN(n694) );
  NOR2_X1 U599 ( .A1(G902), .A2(n355), .ZN(n468) );
  NOR2_X1 U600 ( .A1(G953), .A2(G952), .ZN(n467) );
  NOR2_X1 U601 ( .A1(n468), .A2(n467), .ZN(n469) );
  AND2_X1 U602 ( .A1(n694), .A2(n469), .ZN(n552) );
  INV_X1 U603 ( .A(n476), .ZN(n477) );
  XNOR2_X1 U604 ( .A(KEYINPUT71), .B(n719), .ZN(n516) );
  XOR2_X1 U605 ( .A(n481), .B(n480), .Z(n482) );
  NAND2_X1 U606 ( .A1(n700), .A2(n483), .ZN(n485) );
  NAND2_X1 U607 ( .A1(G210), .A2(n486), .ZN(n484) );
  XNOR2_X2 U608 ( .A(n485), .B(n484), .ZN(n603) );
  INV_X1 U609 ( .A(n603), .ZN(n584) );
  NAND2_X1 U610 ( .A1(G214), .A2(n486), .ZN(n487) );
  XOR2_X1 U611 ( .A(KEYINPUT91), .B(n487), .Z(n681) );
  NAND2_X1 U612 ( .A1(G898), .A2(G953), .ZN(n488) );
  INV_X1 U613 ( .A(n543), .ZN(n530) );
  NAND2_X1 U614 ( .A1(n490), .A2(G221), .ZN(n491) );
  XNOR2_X1 U615 ( .A(n491), .B(KEYINPUT21), .ZN(n668) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n493) );
  XNOR2_X1 U617 ( .A(G140), .B(KEYINPUT96), .ZN(n492) );
  XNOR2_X1 U618 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U619 ( .A(n728), .B(n494), .Z(n497) );
  NAND2_X1 U620 ( .A1(n495), .A2(G214), .ZN(n496) );
  XNOR2_X1 U621 ( .A(n498), .B(KEYINPUT95), .ZN(n502) );
  XNOR2_X1 U622 ( .A(n500), .B(n499), .ZN(n501) );
  NOR2_X1 U623 ( .A1(G902), .A2(n622), .ZN(n505) );
  XNOR2_X1 U624 ( .A(KEYINPUT13), .B(G475), .ZN(n504) );
  NOR2_X1 U625 ( .A1(G902), .A2(n613), .ZN(n507) );
  INV_X1 U626 ( .A(n684), .ZN(n508) );
  INV_X1 U627 ( .A(KEYINPUT65), .ZN(n509) );
  INV_X1 U628 ( .A(n511), .ZN(n512) );
  NAND2_X1 U629 ( .A1(G227), .A2(n355), .ZN(n514) );
  NOR2_X1 U630 ( .A1(G902), .A2(n704), .ZN(n517) );
  INV_X1 U631 ( .A(n590), .ZN(n528) );
  XOR2_X1 U632 ( .A(KEYINPUT81), .B(n528), .Z(n518) );
  NAND2_X1 U633 ( .A1(n518), .A2(n599), .ZN(n519) );
  NOR2_X1 U634 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U635 ( .A(KEYINPUT80), .B(n521), .Z(n522) );
  XNOR2_X1 U636 ( .A(KEYINPUT32), .B(n524), .ZN(n743) );
  NOR2_X1 U637 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U638 ( .A1(n539), .A2(n531), .ZN(n583) );
  INV_X1 U639 ( .A(n740), .ZN(n533) );
  NAND2_X1 U640 ( .A1(n533), .A2(n443), .ZN(n534) );
  NAND2_X1 U641 ( .A1(n535), .A2(n534), .ZN(n548) );
  NOR2_X1 U642 ( .A1(n590), .A2(n669), .ZN(n536) );
  NAND2_X1 U643 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U644 ( .A(KEYINPUT101), .B(n538), .ZN(n742) );
  AND2_X1 U645 ( .A1(n541), .A2(n675), .ZN(n677) );
  NAND2_X1 U646 ( .A1(n677), .A2(n543), .ZN(n542) );
  XNOR2_X1 U647 ( .A(KEYINPUT31), .B(n542), .ZN(n649) );
  NAND2_X1 U648 ( .A1(n561), .A2(n543), .ZN(n544) );
  NOR2_X1 U649 ( .A1(n675), .A2(n544), .ZN(n636) );
  NOR2_X1 U650 ( .A1(n649), .A2(n636), .ZN(n545) );
  NOR2_X1 U651 ( .A1(n686), .A2(n545), .ZN(n546) );
  NOR2_X1 U652 ( .A1(n742), .A2(n546), .ZN(n547) );
  XNOR2_X1 U653 ( .A(KEYINPUT38), .B(n603), .ZN(n682) );
  NAND2_X1 U654 ( .A1(n682), .A2(n681), .ZN(n685) );
  XOR2_X1 U655 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n549) );
  XOR2_X1 U656 ( .A(KEYINPUT108), .B(KEYINPUT28), .Z(n556) );
  NAND2_X1 U657 ( .A1(G953), .A2(G900), .ZN(n551) );
  NAND2_X1 U658 ( .A1(n552), .A2(n551), .ZN(n567) );
  NOR2_X1 U659 ( .A1(n668), .A2(n567), .ZN(n553) );
  XNOR2_X1 U660 ( .A(KEYINPUT70), .B(n553), .ZN(n554) );
  NAND2_X1 U661 ( .A1(n554), .A2(n669), .ZN(n555) );
  NAND2_X1 U662 ( .A1(n558), .A2(n577), .ZN(n559) );
  XOR2_X1 U663 ( .A(KEYINPUT42), .B(n559), .Z(n744) );
  INV_X1 U664 ( .A(KEYINPUT105), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n561), .B(n560), .ZN(n569) );
  NAND2_X1 U666 ( .A1(n562), .A2(n681), .ZN(n565) );
  XOR2_X1 U667 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n563) );
  NAND2_X1 U668 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U669 ( .A1(n586), .A2(n682), .ZN(n573) );
  XNOR2_X1 U670 ( .A(KEYINPUT46), .B(n575), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n577), .A2(n576), .ZN(n644) );
  NOR2_X1 U672 ( .A1(n686), .A2(KEYINPUT47), .ZN(n579) );
  XNOR2_X1 U673 ( .A(n580), .B(KEYINPUT73), .ZN(n582) );
  NAND2_X1 U674 ( .A1(KEYINPUT47), .A2(n644), .ZN(n581) );
  NAND2_X1 U675 ( .A1(n582), .A2(n581), .ZN(n589) );
  NAND2_X1 U676 ( .A1(KEYINPUT47), .A2(n686), .ZN(n587) );
  AND2_X1 U677 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U678 ( .A1(n586), .A2(n585), .ZN(n643) );
  NAND2_X1 U679 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U680 ( .A(KEYINPUT104), .B(n593), .Z(n600) );
  NOR2_X1 U681 ( .A1(n600), .A2(n594), .ZN(n595) );
  NOR2_X1 U682 ( .A1(n596), .A2(n651), .ZN(n597) );
  NOR2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n601), .A2(n681), .ZN(n602) );
  XNOR2_X1 U685 ( .A(n602), .B(KEYINPUT43), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n656) );
  NAND2_X1 U687 ( .A1(n606), .A2(n648), .ZN(n654) );
  NAND2_X1 U688 ( .A1(KEYINPUT2), .A2(n654), .ZN(n607) );
  XNOR2_X1 U689 ( .A(KEYINPUT82), .B(n607), .ZN(n608) );
  NOR2_X1 U690 ( .A1(n611), .A2(n608), .ZN(n609) );
  NAND2_X1 U691 ( .A1(G478), .A2(n707), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT122), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n707), .A2(G217), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(G66) );
  NAND2_X1 U696 ( .A1(n707), .A2(G475), .ZN(n626) );
  XNOR2_X1 U697 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n622), .B(KEYINPUT119), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U701 ( .A(KEYINPUT60), .B(KEYINPUT120), .ZN(n628) );
  XOR2_X1 U702 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n629) );
  XOR2_X1 U703 ( .A(KEYINPUT63), .B(n631), .Z(G57) );
  NAND2_X1 U704 ( .A1(n636), .A2(n387), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(G104), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n634) );
  XNOR2_X1 U707 ( .A(G107), .B(KEYINPUT26), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(n635) );
  XOR2_X1 U709 ( .A(KEYINPUT112), .B(n635), .Z(n638) );
  NAND2_X1 U710 ( .A1(n636), .A2(n648), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G9) );
  XOR2_X1 U712 ( .A(n639), .B(G110), .Z(G12) );
  INV_X1 U713 ( .A(n648), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n640), .A2(n644), .ZN(n642) );
  XNOR2_X1 U715 ( .A(G128), .B(KEYINPUT29), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n642), .B(n641), .ZN(G30) );
  XNOR2_X1 U717 ( .A(G143), .B(n643), .ZN(G45) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U719 ( .A(G146), .B(n646), .Z(G48) );
  NAND2_X1 U720 ( .A1(n649), .A2(n387), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(G113), .ZN(G15) );
  NAND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(G116), .ZN(G18) );
  XNOR2_X1 U724 ( .A(n651), .B(KEYINPUT37), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT114), .ZN(n653) );
  XNOR2_X1 U726 ( .A(G125), .B(n653), .ZN(G27) );
  XOR2_X1 U727 ( .A(G134), .B(n654), .Z(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U729 ( .A(G140), .B(n656), .ZN(G42) );
  NAND2_X1 U730 ( .A1(n712), .A2(n730), .ZN(n658) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n657) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT86), .B(n661), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n680), .A2(n690), .ZN(n662) );
  NOR2_X1 U736 ( .A1(G953), .A2(n662), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n698) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(KEYINPUT50), .B(n667), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n671) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U746 ( .A(KEYINPUT51), .B(n678), .Z(n679) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U754 ( .A(KEYINPUT52), .B(n693), .ZN(n696) );
  NAND2_X1 U755 ( .A1(n694), .A2(G952), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U758 ( .A(KEYINPUT53), .B(n699), .ZN(G75) );
  NAND2_X1 U759 ( .A1(n707), .A2(G210), .ZN(n702) );
  XNOR2_X1 U760 ( .A(n700), .B(n436), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n704), .B(KEYINPUT57), .ZN(n705) );
  XNOR2_X1 U764 ( .A(n706), .B(n705), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U766 ( .A1(n355), .A2(n712), .ZN(n716) );
  NAND2_X1 U767 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U768 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n714), .A2(G898), .ZN(n715) );
  NAND2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n724) );
  XOR2_X1 U771 ( .A(n717), .B(G101), .Z(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n722) );
  NOR2_X1 U773 ( .A1(G898), .A2(n355), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(G69) );
  XOR2_X1 U776 ( .A(n726), .B(n725), .Z(n727) );
  XOR2_X1 U777 ( .A(n728), .B(n727), .Z(n733) );
  INV_X1 U778 ( .A(n733), .ZN(n729) );
  XOR2_X1 U779 ( .A(n729), .B(KEYINPUT124), .Z(n731) );
  XNOR2_X1 U780 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n732), .A2(n355), .ZN(n737) );
  XOR2_X1 U782 ( .A(G227), .B(n733), .Z(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U786 ( .A(G131), .B(KEYINPUT126), .Z(n738) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(G33) );
  XOR2_X1 U788 ( .A(G122), .B(n740), .Z(n741) );
  XNOR2_X1 U789 ( .A(n741), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U790 ( .A(G101), .B(n742), .Z(G3) );
  XOR2_X1 U791 ( .A(n743), .B(G119), .Z(G21) );
  XOR2_X1 U792 ( .A(G137), .B(n744), .Z(G39) );
endmodule

