//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G77), .A2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n203), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n206), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(G250), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n222), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT18), .ZN(new_n250));
  INV_X1    g0050(.A(G169), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n219), .A2(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G87), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n255), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n266), .A2(G232), .A3(new_n253), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT78), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n266), .B1(new_n262), .B2(new_n263), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT78), .ZN(new_n273));
  NOR4_X1   g0073(.A1(new_n272), .A2(new_n273), .A3(new_n269), .A4(new_n255), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n251), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(new_n267), .ZN(new_n276));
  INV_X1    g0076(.A(new_n255), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(new_n270), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n260), .A2(new_n261), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT7), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n226), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT7), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(new_n292), .A3(G68), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n221), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G58), .A2(G68), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G159), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n293), .A2(KEYINPUT16), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n227), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT16), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n283), .A2(new_n226), .A3(KEYINPUT7), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n291), .A2(new_n284), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n294), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n297), .A2(new_n299), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n305), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  OR2_X1    g0111(.A1(KEYINPUT8), .A2(G58), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT8), .A2(G58), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n289), .A2(G1), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n252), .A2(G20), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n303), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n312), .A2(new_n317), .A3(KEYINPUT76), .A4(new_n313), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n314), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(KEYINPUT77), .A3(new_n323), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n304), .A2(new_n310), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n250), .B1(new_n282), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n278), .A2(new_n273), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n268), .A2(KEYINPUT78), .A3(new_n270), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n251), .B1(new_n280), .B2(new_n279), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n326), .A2(new_n327), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n310), .A2(new_n303), .A3(new_n301), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(KEYINPUT18), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(G200), .B1(new_n330), .B2(new_n331), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT79), .B(G190), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n278), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n335), .B(new_n334), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n271), .B2(new_n274), .ZN(new_n347));
  INV_X1    g0147(.A(new_n342), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n328), .A3(KEYINPUT17), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n288), .A2(new_n290), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n257), .A2(G222), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n354), .C1(new_n256), .C2(new_n257), .ZN(new_n355));
  INV_X1    g0155(.A(G77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n283), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(KEYINPUT69), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT69), .B1(new_n355), .B2(new_n357), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n359), .A2(new_n360), .A3(new_n266), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n266), .A2(new_n253), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n277), .B1(new_n362), .B2(new_n219), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT68), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n251), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n226), .A2(G33), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n226), .A2(KEYINPUT70), .A3(G33), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n314), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G150), .ZN(new_n372));
  INV_X1    g0172(.A(new_n298), .ZN(new_n373));
  NOR3_X1   g0173(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(new_n289), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n303), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n303), .A2(new_n315), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G50), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n319), .A2(new_n218), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n360), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n267), .A3(new_n358), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n363), .B(KEYINPUT68), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n280), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n366), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G200), .B1(new_n361), .B2(new_n365), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(new_n383), .A3(G190), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n376), .A2(KEYINPUT9), .A3(new_n378), .A4(new_n379), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT9), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n380), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT10), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n388), .A2(new_n389), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT10), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n392), .A3(new_n396), .A4(new_n387), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n386), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n312), .A2(new_n313), .ZN(new_n399));
  AND2_X1   g0199(.A1(KEYINPUT64), .A2(G20), .ZN(new_n400));
  NOR2_X1   g0200(.A1(KEYINPUT64), .A2(G20), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n399), .A2(new_n298), .B1(new_n402), .B2(G77), .ZN(new_n403));
  OR2_X1    g0203(.A1(KEYINPUT15), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(KEYINPUT15), .A2(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT71), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(KEYINPUT71), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n403), .B1(new_n410), .B2(new_n367), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n303), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n319), .A2(new_n356), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n377), .A2(G77), .ZN(new_n415));
  XOR2_X1   g0215(.A(new_n415), .B(KEYINPUT72), .Z(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT73), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(KEYINPUT73), .A3(new_n412), .A4(new_n413), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G238), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n353), .B(new_n419), .C1(new_n222), .C2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(new_n267), .C1(G107), .C2(new_n353), .ZN(new_n421));
  INV_X1    g0221(.A(new_n362), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G244), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n277), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  INV_X1    g0225(.A(G190), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n418), .B(new_n425), .C1(new_n426), .C2(new_n424), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n352), .B(new_n398), .C1(new_n417), .C2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT75), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  OAI211_X1 g0232(.A(G232), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT74), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n353), .A2(KEYINPUT74), .A3(G232), .A4(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G97), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n353), .A2(G226), .A3(new_n257), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n267), .ZN(new_n440));
  INV_X1    g0240(.A(G238), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n277), .B1(new_n362), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n432), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g0244(.A(KEYINPUT13), .B(new_n442), .C1(new_n439), .C2(new_n267), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n431), .B1(new_n446), .B2(new_n251), .ZN(new_n447));
  OAI221_X1 g0247(.A(G169), .B1(new_n429), .B2(new_n430), .C1(new_n444), .C2(new_n445), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(G179), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n373), .A2(new_n218), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n289), .A2(G68), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n369), .A2(new_n370), .ZN(new_n453));
  AOI211_X1 g0253(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(G77), .ZN(new_n454));
  INV_X1    g0254(.A(new_n303), .ZN(new_n455));
  OR3_X1    g0255(.A1(new_n454), .A2(KEYINPUT11), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT11), .B1(new_n454), .B2(new_n455), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n377), .A2(G68), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n315), .A2(G13), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n460), .A2(KEYINPUT12), .A3(G68), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT12), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n462), .B1(new_n319), .B2(new_n294), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n450), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(G200), .B1(new_n444), .B2(new_n445), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n446), .A2(G190), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n458), .A2(new_n465), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n414), .A2(new_n416), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n424), .A2(new_n251), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(G179), .B2(new_n424), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n467), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n428), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n208), .A2(new_n257), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n210), .A2(G1698), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n477), .B(new_n478), .C1(new_n260), .C2(new_n261), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT86), .A2(G294), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT86), .A2(G294), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(G33), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n267), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  INV_X1    g0285(.A(G45), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(G274), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  NOR2_X1   g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G264), .A3(new_n266), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n484), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT87), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n488), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n426), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n346), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OR3_X1    g0299(.A1(new_n226), .A2(KEYINPUT23), .A3(G107), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n213), .A2(G20), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(KEYINPUT23), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(new_n401), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT64), .A2(G20), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(new_n507), .B1(new_n288), .B2(new_n290), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n508), .B2(G87), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n353), .A2(new_n226), .A3(new_n505), .A4(G87), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n500), .B(new_n504), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(KEYINPUT24), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  INV_X1    g0314(.A(new_n504), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n353), .A2(new_n226), .A3(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n518), .B2(new_n500), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n303), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT25), .B1(new_n319), .B2(new_n213), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n252), .A2(G33), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n455), .A2(new_n460), .A3(new_n524), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n522), .A2(new_n523), .B1(new_n525), .B2(new_n213), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n499), .A2(new_n520), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n512), .A2(KEYINPUT24), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n518), .A2(new_n514), .A3(new_n500), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n455), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n251), .B1(new_n495), .B2(new_n496), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n493), .A2(new_n280), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n531), .A2(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT88), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI221_X1 g0336(.A(KEYINPUT88), .B1(new_n532), .B2(new_n533), .C1(new_n531), .C2(new_n526), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n528), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n353), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n539));
  OAI21_X1  g0339(.A(G244), .B1(new_n260), .B2(new_n261), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n353), .A2(G250), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n257), .B1(new_n545), .B2(KEYINPUT4), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n267), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n491), .A2(new_n266), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G257), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n488), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G200), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n209), .A2(new_n213), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n226), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n373), .A2(new_n356), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n306), .A2(new_n307), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(new_n560), .C1(new_n561), .C2(new_n213), .ZN(new_n562));
  INV_X1    g0362(.A(new_n525), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(new_n303), .B1(G97), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n319), .A2(new_n209), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n547), .A2(G190), .A3(new_n488), .A4(new_n549), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n551), .A2(new_n564), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n550), .A2(new_n251), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(G97), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n213), .B1(new_n306), .B2(new_n307), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n570), .A2(new_n559), .A3(new_n557), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n565), .B(new_n569), .C1(new_n571), .C2(new_n455), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n547), .A2(new_n280), .A3(new_n488), .A4(new_n549), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n353), .A2(KEYINPUT81), .A3(G244), .A4(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n353), .A2(G238), .A3(new_n257), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n501), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n267), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n252), .A2(G45), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n266), .A2(G250), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n266), .A2(KEYINPUT80), .A3(G250), .A4(new_n583), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(G274), .B2(new_n487), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n582), .A2(G179), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n251), .B1(new_n582), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT82), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n582), .A2(G179), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(new_n587), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n487), .A2(G274), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n267), .B2(new_n581), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n592), .B(new_n593), .C1(new_n597), .C2(new_n251), .ZN(new_n598));
  OAI211_X1 g0398(.A(G33), .B(G97), .C1(new_n400), .C2(new_n401), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n400), .A2(new_n401), .B1(new_n600), .B2(new_n437), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n554), .A2(new_n207), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n353), .A2(new_n226), .A3(G68), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n303), .ZN(new_n607));
  INV_X1    g0407(.A(new_n410), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n563), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n410), .A2(new_n319), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT83), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n606), .A2(new_n303), .B1(new_n319), .B2(new_n410), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n609), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n591), .A2(new_n598), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n582), .A2(new_n588), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n582), .A2(G190), .A3(new_n588), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n563), .A2(G87), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n613), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(KEYINPUT85), .A2(KEYINPUT21), .ZN(new_n624));
  INV_X1    g0424(.A(G116), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n319), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n455), .A2(new_n460), .A3(G116), .A4(new_n524), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n287), .A2(G97), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n628), .B(new_n543), .C1(new_n400), .C2(new_n401), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n302), .A2(new_n227), .B1(G20), .B2(new_n625), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n629), .A2(KEYINPUT20), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT20), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n626), .B(new_n627), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT84), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n548), .A2(G270), .ZN(new_n635));
  INV_X1    g0435(.A(G303), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n266), .B1(new_n283), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n353), .B1(new_n214), .B2(new_n257), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n210), .A2(G1698), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n635), .A2(new_n640), .A3(new_n488), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G169), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n624), .B1(new_n634), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n642), .ZN(new_n644));
  INV_X1    g0444(.A(new_n624), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT84), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n633), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n633), .A2(new_n646), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n644), .B(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n641), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n651), .B(G179), .C1(new_n648), .C2(new_n649), .ZN(new_n652));
  INV_X1    g0452(.A(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n341), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n641), .A2(G200), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n647), .A4(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n643), .A2(new_n650), .A3(new_n652), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n623), .A2(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n476), .A2(new_n538), .A3(new_n575), .A4(new_n658), .ZN(G372));
  AND3_X1   g0459(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n613), .A2(new_n614), .A3(new_n609), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n614), .B1(new_n613), .B2(new_n609), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n662), .A2(new_n663), .B1(new_n589), .B2(new_n590), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n660), .A2(new_n661), .A3(new_n622), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n617), .A2(new_n660), .A3(new_n622), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(KEYINPUT26), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n531), .A2(new_n526), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n499), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n613), .A2(new_n621), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(G200), .B2(new_n618), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n593), .B1(new_n597), .B2(new_n251), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n620), .A2(new_n672), .B1(new_n616), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n575), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n534), .A2(new_n643), .A3(new_n650), .A4(new_n652), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT89), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n567), .A2(new_n664), .A3(new_n574), .A4(new_n622), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n528), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n534), .A2(new_n643), .A3(new_n650), .A4(new_n652), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n668), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n476), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n394), .A2(new_n397), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT90), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n338), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n329), .A2(new_n337), .A3(KEYINPUT90), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n471), .A2(new_n473), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n470), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n351), .B1(new_n692), .B2(new_n467), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n685), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(new_n385), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT91), .ZN(G369));
  NOR2_X1   g0497(.A1(new_n402), .A2(new_n318), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .A3(G1), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT27), .B1(new_n699), .B2(G1), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(G213), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n634), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n657), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n643), .A2(new_n650), .A3(new_n652), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n706), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n538), .B1(new_n669), .B2(new_n705), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n534), .B2(new_n705), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n534), .A2(new_n704), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n708), .A2(new_n705), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n717), .B1(new_n719), .B2(new_n538), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n204), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n603), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n229), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT89), .B1(new_n675), .B2(new_n676), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n680), .A2(new_n678), .A3(new_n681), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n704), .B1(new_n731), .B2(new_n668), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n593), .A2(new_n493), .ZN(new_n735));
  INV_X1    g0535(.A(new_n550), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n635), .A2(new_n640), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n493), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n582), .B2(new_n588), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n280), .A3(new_n550), .A4(new_n641), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n739), .A2(new_n582), .A3(G179), .A4(new_n588), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n737), .A2(new_n547), .A3(new_n488), .A4(new_n549), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n738), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT31), .B1(new_n746), .B2(new_n704), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(KEYINPUT92), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT92), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(new_n747), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n658), .A2(new_n538), .A3(new_n575), .A4(new_n705), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT29), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n664), .A2(new_n622), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT26), .B1(new_n759), .B2(new_n574), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n617), .A2(new_n661), .A3(new_n660), .A4(new_n622), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(new_n761), .A3(new_n664), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n536), .A2(new_n537), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n680), .B1(new_n764), .B2(new_n708), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT93), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n760), .A2(new_n761), .A3(new_n766), .A4(new_n664), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n763), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n758), .B1(new_n768), .B2(new_n705), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n734), .A2(new_n757), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n728), .B1(new_n770), .B2(G1), .ZN(G364));
  AOI21_X1  g0571(.A(new_n227), .B1(G20), .B2(new_n251), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n226), .A2(new_n280), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G200), .A3(new_n341), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  INV_X1    g0576(.A(G326), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n774), .A2(new_n426), .A3(new_n346), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n774), .A2(new_n346), .A3(new_n341), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT95), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n774), .A2(KEYINPUT95), .A3(new_n346), .A4(new_n341), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n402), .A2(new_n426), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT97), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(G179), .A3(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G329), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n791), .A2(G179), .A3(new_n346), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n774), .A2(new_n426), .A3(G200), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  OAI21_X1  g0599(.A(new_n283), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n780), .A2(new_n788), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n346), .A2(G179), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G20), .A3(G190), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n480), .A2(new_n481), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n426), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n226), .A2(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n801), .B1(new_n636), .B2(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT99), .Z(new_n808));
  INV_X1    g0608(.A(new_n775), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n283), .B1(new_n809), .B2(G50), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n207), .B2(new_n803), .C1(new_n213), .C2(new_n795), .ZN(new_n811));
  INV_X1    g0611(.A(new_n806), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G97), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n779), .B2(new_n356), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n792), .ZN(new_n816));
  INV_X1    g0616(.A(G159), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT32), .ZN(new_n819));
  INV_X1    g0619(.A(new_n798), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n818), .A2(new_n819), .B1(G68), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n815), .B(new_n821), .C1(new_n819), .C2(new_n818), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n785), .B(KEYINPUT96), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(G58), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n772), .B1(new_n808), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n698), .A2(G45), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(new_n724), .A3(G1), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT100), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n711), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n353), .A2(G355), .A3(new_n204), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n245), .A2(new_n486), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n722), .A2(new_n353), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G45), .B2(new_n229), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n834), .B1(G116), .B2(new_n204), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n831), .A2(new_n772), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n825), .A2(new_n828), .A3(new_n833), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n710), .A2(G330), .ZN(new_n842));
  OR3_X1    g0642(.A1(new_n713), .A2(new_n828), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(G396));
  INV_X1    g0644(.A(new_n772), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n294), .A2(new_n795), .B1(new_n816), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n823), .A2(G143), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n809), .B1(new_n820), .B2(G150), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n817), .C2(new_n779), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n851));
  AOI211_X1 g0651(.A(new_n283), .B(new_n847), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n803), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(G50), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n855), .B1(new_n221), .B2(new_n806), .C1(new_n851), .C2(new_n850), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n809), .A2(G303), .B1(G97), .B2(new_n812), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n857), .B1(new_n213), .B2(new_n803), .C1(new_n796), .C2(new_n798), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n785), .A2(G294), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n795), .A2(new_n207), .ZN(new_n860));
  NOR4_X1   g0660(.A1(new_n858), .A2(new_n353), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n625), .B2(new_n779), .C1(new_n778), .C2(new_n816), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT101), .Z(new_n863));
  AOI21_X1  g0663(.A(new_n845), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n414), .A2(new_n416), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n704), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n427), .B2(new_n417), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n474), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n691), .A2(new_n705), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n830), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n864), .A2(new_n827), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n772), .A2(new_n829), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(G77), .B2(new_n875), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n704), .B(new_n870), .C1(new_n731), .C2(new_n668), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT103), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n870), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n877), .B1(new_n733), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n757), .B1(new_n880), .B2(KEYINPUT104), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n880), .B(KEYINPUT104), .Z(new_n882));
  OAI211_X1 g0682(.A(new_n827), .B(new_n881), .C1(new_n882), .C2(new_n757), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n883), .ZN(G384));
  OAI21_X1  g0684(.A(new_n476), .B1(new_n734), .B2(new_n769), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n695), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n466), .A2(new_n704), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n467), .A2(new_n887), .A3(new_n470), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n450), .A2(new_n466), .A3(new_n704), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n683), .A2(new_n705), .A3(new_n871), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n869), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT106), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n336), .A2(new_n895), .A3(new_n275), .A4(new_n281), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  INV_X1    g0697(.A(new_n702), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n336), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n343), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n895), .B1(new_n333), .B2(new_n336), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n336), .B1(new_n347), .B2(new_n348), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n293), .B2(new_n300), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n324), .B1(new_n304), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n282), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n903), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n343), .B(KEYINPUT105), .C1(new_n282), .C2(new_n907), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n907), .A2(new_n702), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n902), .B1(new_n913), .B2(KEYINPUT37), .ZN(new_n914));
  INV_X1    g0714(.A(new_n351), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n915), .B2(new_n338), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n894), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n911), .B1(new_n339), .B2(new_n351), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n301), .A2(new_n303), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n323), .B(new_n322), .C1(new_n919), .C2(new_n905), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n333), .A2(new_n920), .B1(new_n349), .B2(new_n328), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n911), .B1(new_n921), .B2(KEYINPUT105), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n897), .B1(new_n922), .B2(new_n909), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT38), .B(new_n918), .C1(new_n923), .C2(new_n902), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n893), .A2(new_n925), .ZN(new_n926));
  AND4_X1   g0726(.A1(new_n897), .A2(new_n896), .A3(new_n343), .A4(new_n899), .ZN(new_n927));
  INV_X1    g0727(.A(new_n901), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n343), .B(new_n899), .C1(new_n328), .C2(new_n282), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n927), .A2(new_n928), .B1(KEYINPUT37), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n329), .A2(new_n337), .A3(KEYINPUT90), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT90), .B1(new_n329), .B2(new_n337), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n915), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n899), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n924), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n467), .A2(new_n704), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n924), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n690), .A2(new_n702), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n926), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n886), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n752), .A2(new_n747), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n754), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n870), .B1(new_n888), .B2(new_n889), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n925), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n947), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n899), .B1(new_n689), .B2(new_n915), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n894), .B1(new_n952), .B2(new_n930), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n953), .B2(new_n924), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n954), .B2(new_n949), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n955), .A2(new_n946), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n949), .B1(new_n936), .B2(new_n948), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n924), .B2(new_n917), .ZN(new_n959));
  OAI21_X1  g0759(.A(G330), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n712), .B1(new_n754), .B2(new_n945), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n476), .A2(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n956), .A2(new_n476), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n944), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n252), .B2(new_n698), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n555), .A2(new_n556), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n625), .B1(new_n966), .B2(KEYINPUT35), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n228), .C1(KEYINPUT35), .C2(new_n966), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT36), .ZN(new_n969));
  OAI21_X1  g0769(.A(G77), .B1(new_n221), .B2(new_n294), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n970), .A2(new_n229), .B1(G50), .B2(new_n294), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(G1), .A3(new_n318), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n965), .A2(new_n969), .A3(new_n972), .ZN(G367));
  NAND2_X1  g0773(.A1(new_n704), .A2(new_n572), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n575), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n660), .A2(new_n704), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n719), .A2(new_n538), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n536), .A2(new_n537), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n574), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n705), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT108), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n704), .A2(new_n671), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n759), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n616), .A3(new_n673), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  INV_X1    g0791(.A(new_n990), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n986), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n986), .A2(new_n995), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n716), .B2(new_n978), .ZN(new_n999));
  INV_X1    g0799(.A(new_n716), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n1000), .A3(new_n977), .A4(new_n997), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n723), .B(KEYINPUT41), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n715), .A2(new_n719), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT110), .B2(new_n979), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT110), .B2(new_n979), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n713), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n720), .A2(new_n977), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n720), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT44), .B1(new_n720), .B2(new_n977), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1009), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1011), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1014), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1008), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1007), .A2(new_n770), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1003), .B1(new_n1019), .B2(new_n770), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n826), .A2(G1), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT111), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n999), .B(new_n1001), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n836), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n839), .B1(new_n204), .B2(new_n410), .C1(new_n235), .C2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n827), .B1(new_n992), .B2(new_n832), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n776), .A2(new_n778), .B1(new_n796), .B2(new_n779), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n804), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n820), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n823), .A2(G303), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n792), .A2(G317), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n794), .A2(G97), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n213), .B2(new_n806), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT46), .B1(new_n803), .B2(new_n625), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n803), .A2(KEYINPUT46), .A3(new_n625), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n353), .B(new_n1034), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n795), .A2(new_n356), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n353), .B1(new_n221), .B2(new_n803), .C1(new_n779), .C2(new_n218), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G137), .C2(new_n792), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n812), .A2(G68), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n776), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1043), .A2(G143), .B1(G159), .B2(new_n820), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n785), .A2(G150), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT47), .Z(new_n1048));
  OAI211_X1 g0848(.A(new_n1026), .B(new_n1027), .C1(new_n1048), .C2(new_n845), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1024), .A2(new_n1049), .ZN(G387));
  AOI22_X1  g0850(.A1(new_n823), .A2(G317), .B1(G311), .B2(new_n820), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n636), .B2(new_n779), .C1(new_n787), .C2(new_n776), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT48), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n812), .A2(G283), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n853), .A2(new_n1029), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n283), .B1(new_n816), .B2(new_n777), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G116), .B2(new_n794), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n608), .A2(new_n812), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n786), .B2(new_n218), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT113), .Z(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G159), .B2(new_n809), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n283), .B1(new_n853), .B2(G77), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1033), .B(new_n1068), .C1(new_n816), .C2(new_n372), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT112), .Z(new_n1070));
  INV_X1    g0870(.A(new_n779), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(G68), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n820), .A2(new_n399), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n845), .B1(new_n1063), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n314), .A2(G50), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(G68), .A2(G77), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1077), .A2(new_n486), .A3(new_n1078), .A4(new_n725), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1025), .B1(new_n240), .B2(G45), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n725), .A2(new_n283), .A3(new_n722), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n722), .A2(new_n213), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n772), .B(new_n831), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n832), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n715), .A2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1075), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(new_n828), .B1(new_n1007), .B2(new_n1023), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1007), .A2(new_n770), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1007), .A2(new_n770), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n723), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(G393));
  NOR2_X1   g0892(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(new_n716), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n723), .A3(new_n1019), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1094), .A2(new_n1022), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n839), .B1(new_n209), .B2(new_n204), .C1(new_n248), .C2(new_n1025), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n977), .A2(G20), .A3(new_n830), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n785), .A2(G159), .B1(G150), .B2(new_n809), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n806), .A2(new_n356), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n860), .B1(G143), .B2(new_n792), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n353), .C1(new_n294), .C2(new_n803), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n218), .B2(new_n798), .C1(new_n314), .C2(new_n779), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n816), .A2(new_n787), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n785), .A2(G311), .B1(G317), .B2(new_n809), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT52), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(new_n353), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1071), .A2(G294), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n820), .A2(G303), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n795), .A2(new_n213), .B1(new_n796), .B2(new_n803), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G116), .B2(new_n812), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1109), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n827), .B(new_n1099), .C1(new_n1118), .C2(new_n772), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1097), .B1(new_n1098), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1096), .A2(new_n1120), .ZN(G390));
  NAND2_X1  g0921(.A1(new_n938), .A2(new_n940), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n829), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n874), .A2(new_n314), .ZN(new_n1124));
  INV_X1    g0924(.A(G137), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n353), .B1(new_n798), .B2(new_n1125), .C1(new_n795), .C2(new_n218), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT54), .B(G143), .Z(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1071), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n785), .A2(G132), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n803), .A2(new_n372), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n775), .A2(new_n1132), .B1(new_n817), .B2(new_n806), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G125), .B2(new_n792), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n798), .A2(new_n213), .B1(new_n207), .B2(new_n803), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1102), .B(new_n1136), .C1(G283), .C2(new_n809), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n792), .A2(G294), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n785), .A2(G116), .B1(G68), .B2(new_n794), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n283), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n779), .A2(new_n209), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT120), .Z(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n772), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1123), .A2(new_n828), .A3(new_n1124), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT39), .B1(new_n953), .B2(new_n924), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n924), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n893), .A2(new_n939), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n768), .A2(new_n705), .A3(new_n868), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n869), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n890), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n939), .B1(new_n953), .B2(new_n924), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n755), .A2(G330), .A3(new_n947), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1148), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n732), .A2(new_n868), .B1(new_n691), .B2(new_n705), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1156), .A2(new_n891), .B1(new_n467), .B2(new_n704), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1157), .A2(new_n1122), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n961), .A2(new_n947), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1145), .B1(new_n1160), .B2(new_n1022), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT121), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT117), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n879), .B1(new_n1164), .B2(new_n961), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n946), .A2(G330), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT117), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n890), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1154), .A2(new_n1149), .A3(new_n869), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT118), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n870), .B(KEYINPUT103), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1166), .B2(KEYINPUT117), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n961), .A2(new_n1164), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n891), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT118), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1154), .A2(new_n869), .A3(new_n1149), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n891), .B1(new_n756), .B2(new_n870), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1159), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1156), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT116), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n962), .B(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n885), .A3(new_n695), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT119), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1148), .A2(new_n1154), .A3(new_n1153), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1159), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1188), .A2(KEYINPUT119), .A3(new_n1160), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n723), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1163), .A2(new_n1195), .ZN(G378));
  AOI21_X1  g0996(.A(new_n1186), .B1(new_n1192), .B2(new_n1183), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n685), .A2(new_n385), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1199), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n398), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1200), .A2(new_n380), .A3(new_n898), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n898), .A2(new_n380), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n398), .A2(new_n1201), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1199), .B(new_n386), .C1(new_n394), .C2(new_n397), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n960), .A2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1203), .A2(new_n1207), .A3(KEYINPUT122), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT122), .B1(new_n1203), .B2(new_n1207), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(G330), .C1(new_n957), .C2(new_n959), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1210), .A2(new_n943), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n943), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n723), .B1(new_n1197), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT124), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1170), .A2(new_n1177), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1187), .B1(new_n1160), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT123), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n943), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1214), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1208), .B1(new_n955), .B2(G330), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1210), .A2(new_n943), .A3(new_n1214), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1222), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1216), .A2(KEYINPUT123), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1221), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT124), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(new_n723), .C1(new_n1197), .C2(new_n1217), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1219), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n786), .A2(new_n213), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G41), .B1(new_n1071), .B2(new_n608), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n812), .A2(G68), .B1(G77), .B2(new_n853), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n625), .C2(new_n775), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n795), .A2(new_n221), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1236), .A2(new_n1239), .A3(new_n353), .A4(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n209), .B2(new_n798), .C1(new_n796), .C2(new_n816), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT58), .Z(new_n1243));
  OAI21_X1  g1043(.A(new_n218), .B1(new_n260), .B2(G41), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n798), .A2(new_n846), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n812), .A2(G150), .B1(new_n853), .B2(new_n1127), .ZN(new_n1246));
  INV_X1    g1046(.A(G125), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1246), .B1(new_n775), .B2(new_n1247), .C1(new_n1125), .C2(new_n779), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1245), .B(new_n1248), .C1(G128), .C2(new_n785), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT59), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G33), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G41), .B1(new_n792), .B2(G124), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n817), .C2(new_n795), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1244), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n772), .B1(new_n1243), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n874), .A2(new_n218), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1213), .A2(new_n829), .ZN(new_n1258));
  AND4_X1   g1058(.A1(new_n828), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1260), .B2(new_n1023), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1235), .A2(new_n1261), .ZN(G375));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1022), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n816), .A2(new_n1132), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n823), .A2(G137), .B1(new_n820), .B2(new_n1127), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n353), .B1(new_n779), .B2(new_n372), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1267), .B(new_n1240), .C1(G132), .C2(new_n809), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(new_n218), .C2(new_n806), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1265), .B(new_n1269), .C1(G159), .C2(new_n853), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1064), .B1(new_n209), .B2(new_n803), .C1(new_n779), .C2(new_n213), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n353), .B(new_n1271), .C1(G116), .C2(new_n820), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1039), .B1(new_n785), .B2(G283), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1272), .B(new_n1273), .C1(new_n636), .C2(new_n816), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G294), .B2(new_n809), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n772), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n874), .A2(new_n294), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n891), .A2(new_n829), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1276), .A2(new_n828), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1263), .B1(new_n1264), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(KEYINPUT125), .B(new_n1279), .C1(new_n1220), .C2(new_n1022), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1003), .B1(new_n1220), .B2(new_n1186), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1188), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(G381));
  INV_X1    g1086(.A(new_n1161), .ZN(new_n1287));
  AND4_X1   g1087(.A1(new_n1195), .A2(new_n1235), .A3(new_n1287), .A4(new_n1261), .ZN(new_n1288));
  INV_X1    g1088(.A(G384), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1024), .A2(new_n1049), .A3(new_n1120), .A4(new_n1096), .ZN(new_n1291));
  INV_X1    g1091(.A(G396), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1088), .A2(new_n1292), .A3(new_n1091), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(KEYINPUT126), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1290), .A2(new_n1294), .A3(new_n1297), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1296), .A2(new_n1298), .ZN(G407));
  NAND2_X1  g1099(.A1(new_n1288), .A2(new_n703), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G213), .B(new_n1300), .C1(new_n1296), .C2(new_n1298), .ZN(G409));
  INV_X1    g1101(.A(KEYINPUT60), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1220), .A2(KEYINPUT60), .A3(new_n1186), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1188), .A3(new_n723), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1283), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1289), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1283), .A2(new_n1305), .A3(G384), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n703), .A2(G213), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1309), .A2(KEYINPUT127), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1307), .A2(new_n1308), .A3(new_n1313), .A4(new_n1310), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1235), .A2(G378), .A3(new_n1261), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1259), .B1(new_n1320), .B2(new_n1023), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1321), .B1(new_n1230), .B2(new_n1003), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1195), .A3(new_n1287), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1309), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1325), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G393), .A2(G396), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1293), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G387), .A2(G390), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1291), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1291), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1312), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1328), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1336), .A2(KEYINPUT63), .A3(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1326), .A2(new_n1329), .A3(new_n1335), .A4(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT62), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1336), .A2(new_n1340), .A3(new_n1337), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1342), .B1(new_n1336), .B2(new_n1317), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1340), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1339), .B1(new_n1345), .B2(new_n1335), .ZN(G405));
  NAND3_X1  g1146(.A1(G375), .A2(new_n1195), .A3(new_n1287), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1319), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1337), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1347), .A2(new_n1328), .A3(new_n1319), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  OR2_X1    g1151(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1351), .B(new_n1352), .ZN(G402));
endmodule


