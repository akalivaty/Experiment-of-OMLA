//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n212), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(G77), .Z(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n214), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n217), .B(new_n221), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n231), .A2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G169), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n259), .A3(G226), .ZN(new_n260));
  INV_X1    g0060(.A(G232), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n255), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G97), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT76), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT76), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT69), .B(G1698), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n262), .B1(new_n269), .B2(G226), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n268), .B(new_n265), .C1(new_n270), .C2(new_n255), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n277), .A3(G274), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(G238), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n273), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n252), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT14), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n273), .A2(new_n285), .A3(new_n282), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n273), .B2(new_n282), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n287), .A2(new_n288), .B1(new_n291), .B2(G179), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT78), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n287), .B2(new_n288), .ZN(new_n294));
  OAI211_X1 g0094(.A(KEYINPUT78), .B(KEYINPUT14), .C1(new_n291), .C2(new_n252), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n219), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n211), .B2(G20), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G68), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT77), .ZN(new_n301));
  INV_X1    g0101(.A(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n212), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT72), .B1(G20), .B2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G50), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n304), .A2(G20), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G13), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n314), .A2(new_n212), .A3(G1), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n202), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT12), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(KEYINPUT11), .B2(new_n311), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n291), .A2(G190), .ZN(new_n322));
  OAI21_X1  g0122(.A(G200), .B1(new_n289), .B2(new_n290), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(new_n269), .A3(G222), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(G1698), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT70), .B(G223), .Z(new_n331));
  OAI221_X1 g0131(.A(new_n329), .B1(new_n222), .B2(new_n328), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n272), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n279), .B1(G226), .B2(new_n281), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(G200), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT10), .ZN(new_n340));
  INV_X1    g0140(.A(new_n315), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(G50), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n299), .B2(G50), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n208), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n307), .A2(G150), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n212), .A2(G33), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT8), .B(G58), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT8), .ZN(new_n350));
  OR3_X1    g0150(.A1(new_n350), .A2(KEYINPUT71), .A3(G58), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n344), .B1(new_n353), .B2(new_n298), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n339), .A2(new_n340), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n337), .A2(new_n357), .A3(new_n338), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT10), .B1(new_n359), .B2(new_n355), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n353), .A2(new_n298), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n343), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n364), .C1(new_n336), .C2(G169), .ZN(new_n365));
  AOI21_X1  g0165(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT73), .B1(new_n354), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT74), .B(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n336), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT75), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT75), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n299), .A2(G77), .ZN(new_n375));
  INV_X1    g0175(.A(new_n222), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n341), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n376), .A2(G20), .B1(new_n379), .B2(new_n309), .ZN(new_n380));
  INV_X1    g0180(.A(new_n348), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n307), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n298), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n255), .A2(G107), .ZN(new_n385));
  OAI21_X1  g0185(.A(G238), .B1(new_n253), .B2(new_n254), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n257), .B(new_n259), .C1(new_n253), .C2(new_n254), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n385), .B1(new_n386), .B2(new_n256), .C1(new_n261), .C2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n388), .A2(new_n272), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n278), .B1(new_n280), .B2(new_n223), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n384), .B1(new_n392), .B2(new_n252), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n368), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(G190), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n384), .C1(new_n397), .C2(new_n391), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n361), .A2(new_n374), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n326), .A2(new_n212), .A3(new_n327), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n202), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n203), .A2(new_n205), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G20), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n307), .A2(G159), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n401), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n255), .B2(new_n212), .ZN(new_n413));
  NOR4_X1   g0213(.A1(new_n253), .A2(new_n254), .A3(new_n403), .A4(G20), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n408), .A2(G20), .B1(new_n307), .B2(G159), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(KEYINPUT16), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n417), .A3(new_n298), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n352), .A2(new_n341), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n299), .B2(new_n352), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n278), .B1(new_n280), .B2(new_n261), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G226), .A2(G1698), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n269), .B2(G223), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n423), .B1(new_n426), .B2(new_n255), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n427), .B2(new_n272), .ZN(new_n428));
  INV_X1    g0228(.A(new_n368), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n257), .A2(new_n259), .A3(G223), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n255), .B1(new_n431), .B2(new_n424), .ZN(new_n432));
  INV_X1    g0232(.A(new_n423), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n272), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G274), .ZN(new_n435));
  INV_X1    g0235(.A(new_n219), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n276), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n281), .A2(G232), .B1(new_n437), .B2(new_n275), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n421), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n420), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n415), .A2(new_n416), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n302), .B1(new_n449), .B2(new_n401), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(new_n417), .ZN(new_n451));
  INV_X1    g0251(.A(G190), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n434), .A2(new_n452), .A3(new_n438), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n428), .B2(G200), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(KEYINPUT17), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n418), .A3(new_n420), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT18), .B1(new_n421), .B2(new_n441), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT79), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n447), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n325), .A2(new_n400), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n379), .A2(new_n341), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n211), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n341), .A2(new_n302), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G87), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR3_X1   g0272(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(G20), .B1(G33), .B2(G97), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT19), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n309), .A2(new_n476), .A3(G97), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(new_n326), .B2(new_n327), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n475), .A2(new_n477), .B1(new_n478), .B2(G68), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n298), .B1(new_n479), .B2(KEYINPUT83), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n328), .A2(new_n212), .A3(G68), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G97), .A2(G107), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n470), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n265), .A2(new_n212), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n347), .A2(KEYINPUT19), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n481), .B(KEYINPUT83), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n467), .B(new_n472), .C1(new_n480), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n211), .A2(G45), .ZN(new_n491));
  INV_X1    g0291(.A(G250), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n211), .A2(new_n435), .A3(G45), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n277), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n257), .A2(new_n259), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n386), .C2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n500), .B2(new_n272), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n397), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n465), .B1(new_n490), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n481), .B1(new_n485), .B2(new_n487), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n302), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n466), .B1(new_n506), .B2(new_n488), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(new_n272), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n495), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n507), .A2(KEYINPUT84), .A3(new_n510), .A4(new_n472), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(G190), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n503), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n387), .B2(new_n223), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n328), .A2(new_n269), .A3(KEYINPUT4), .A4(G244), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G283), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G250), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n328), .A2(KEYINPUT81), .A3(G250), .A4(G1698), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n272), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT5), .B(G41), .ZN(new_n525));
  INV_X1    g0325(.A(new_n491), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(new_n436), .B2(new_n276), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G257), .ZN(new_n528));
  OR2_X1    g0328(.A1(KEYINPUT5), .A2(G41), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT5), .A2(G41), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n491), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n437), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n524), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n521), .A2(new_n522), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(new_n516), .A3(new_n517), .A4(new_n515), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n533), .B1(new_n538), .B2(new_n272), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G190), .ZN(new_n540));
  OAI21_X1  g0340(.A(G107), .B1(new_n413), .B2(new_n414), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  AND2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n482), .ZN(new_n544));
  INV_X1    g0344(.A(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n307), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n302), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n341), .A2(G97), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n469), .B2(new_n486), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT80), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n307), .A2(G77), .ZN(new_n554));
  INV_X1    g0354(.A(new_n546), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n542), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n554), .B1(new_n557), .B2(new_n212), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n545), .B1(new_n404), .B2(new_n405), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n298), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT80), .ZN(new_n561));
  INV_X1    g0361(.A(new_n469), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n550), .B1(new_n562), .B2(G97), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n536), .A2(new_n540), .A3(new_n553), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n501), .A2(new_n368), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI221_X1 g0368(.A(new_n467), .B1(new_n378), .B2(new_n469), .C1(new_n480), .C2(new_n489), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n501), .A2(new_n368), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n501), .A2(G169), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n568), .B(new_n569), .C1(new_n572), .C2(new_n567), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n368), .B(new_n533), .C1(new_n538), .C2(new_n272), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n252), .B1(new_n524), .B2(new_n534), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n574), .A2(new_n575), .B1(new_n549), .B2(new_n552), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n513), .A2(new_n565), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n212), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n328), .A2(new_n580), .A3(new_n212), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n498), .A2(G20), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n212), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n545), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n583), .B1(new_n582), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n298), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT25), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n545), .B1(new_n592), .B2(KEYINPUT25), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n341), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n315), .A2(new_n592), .A3(KEYINPUT25), .A4(new_n545), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n562), .A2(G107), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G294), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n599), .B(new_n600), .C1(new_n387), .C2(new_n492), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n272), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n527), .A2(G264), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n532), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(KEYINPUT87), .A3(G169), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n601), .A2(new_n272), .B1(G264), .B2(new_n527), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G179), .A3(new_n532), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT87), .B1(new_n604), .B2(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n598), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n604), .A2(G190), .ZN(new_n611));
  AOI21_X1  g0411(.A(G200), .B1(new_n606), .B2(new_n532), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n591), .B(new_n597), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT88), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT88), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n326), .A2(G303), .A3(new_n327), .ZN(new_n619));
  OAI21_X1  g0419(.A(G257), .B1(new_n253), .B2(new_n254), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n499), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n272), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n527), .A2(G270), .B1(new_n437), .B2(new_n531), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(KEYINPUT21), .A3(G169), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(G179), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n341), .A2(G116), .A3(new_n302), .A4(new_n468), .ZN(new_n628));
  INV_X1    g0428(.A(G116), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n315), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n297), .A2(new_n219), .B1(G20), .B2(new_n629), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n517), .B(new_n212), .C1(G33), .C2(new_n486), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n631), .A2(KEYINPUT20), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT20), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n628), .B(new_n630), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n624), .B2(G200), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n452), .B2(new_n624), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n624), .A2(G169), .A3(new_n635), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT85), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n636), .B(new_n638), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n615), .A2(new_n617), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n464), .A2(new_n577), .A3(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n395), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n296), .A2(new_n320), .B1(new_n324), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n455), .A2(new_n458), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n648), .A2(new_n649), .B1(new_n460), .B2(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n361), .B1(new_n372), .B2(new_n373), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n572), .A2(new_n569), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AOI211_X1 g0454(.A(new_n466), .B(new_n471), .C1(new_n506), .C2(new_n488), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT89), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n509), .A2(new_n656), .A3(G200), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT89), .B1(new_n501), .B2(new_n397), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n655), .A2(new_n512), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n613), .A3(new_n653), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n639), .A2(new_n640), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT85), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n640), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n627), .B2(new_n635), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n660), .B1(new_n610), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n565), .A2(new_n576), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n654), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n657), .A2(new_n512), .A3(new_n658), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n469), .A2(new_n378), .ZN(new_n671));
  AOI211_X1 g0471(.A(new_n671), .B(new_n466), .C1(new_n506), .C2(new_n488), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n566), .B1(G169), .B2(new_n501), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n670), .A2(new_n490), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n549), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n561), .B1(new_n560), .B2(new_n563), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n574), .A2(new_n575), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n669), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n535), .A2(G169), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n539), .A2(new_n429), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n553), .A2(new_n564), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n659), .A2(new_n682), .A3(new_n683), .A4(new_n653), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT90), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n669), .ZN(new_n686));
  INV_X1    g0486(.A(new_n576), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(KEYINPUT26), .A3(new_n573), .A4(new_n513), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n679), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n668), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n652), .B1(new_n464), .B2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n635), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n644), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n635), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT91), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(new_n707), .A3(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n610), .A2(new_n616), .A3(new_n613), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n616), .B1(new_n610), .B2(new_n613), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n598), .A2(new_n698), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n610), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n698), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n698), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n701), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n710), .A2(new_n720), .A3(new_n711), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n715), .B2(new_n719), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(G399));
  INV_X1    g0523(.A(new_n215), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G41), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n483), .A2(G116), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G1), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n218), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(new_n726), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT92), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n565), .A2(new_n576), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT95), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n665), .A2(new_n610), .ZN(new_n737));
  INV_X1    g0537(.A(new_n660), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n565), .A2(new_n576), .A3(KEYINPUT95), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n513), .A2(new_n573), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n669), .A3(new_n687), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n654), .B1(new_n684), .B2(KEYINPUT26), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n733), .B1(new_n744), .B2(new_n719), .ZN(new_n745));
  AOI211_X1 g0545(.A(KEYINPUT29), .B(new_n698), .C1(new_n668), .C2(new_n689), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n577), .A2(new_n698), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n712), .A2(new_n747), .A3(new_n644), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n606), .A2(new_n501), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n622), .A2(new_n623), .A3(G179), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n539), .A2(new_n749), .A3(KEYINPUT30), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT93), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n606), .A2(new_n501), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n626), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(KEYINPUT93), .A3(KEYINPUT30), .A4(new_n539), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(new_n501), .A3(new_n606), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(new_n535), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n501), .A2(new_n429), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n535), .A2(new_n604), .A3(new_n624), .A4(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n753), .A2(new_n756), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(KEYINPUT94), .A3(KEYINPUT31), .A4(new_n698), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n698), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT94), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n748), .A2(new_n763), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n745), .B(new_n746), .C1(G330), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n732), .B1(new_n771), .B2(G1), .ZN(G364));
  NOR2_X1   g0572(.A1(new_n314), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n211), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n725), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n704), .B2(new_n705), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n708), .A3(new_n706), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n776), .B(KEYINPUT96), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n724), .A2(new_n255), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G355), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G116), .B2(new_n215), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n724), .A2(new_n328), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT97), .Z(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G45), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(new_n218), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n247), .A2(new_n786), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n219), .B1(G20), .B2(new_n252), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n779), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n793), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n368), .A2(new_n212), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT99), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n368), .A2(KEYINPUT99), .A3(new_n212), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n452), .B(new_n397), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(G190), .B(new_n397), .C1(new_n800), .C2(new_n801), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G311), .A2(new_n803), .B1(new_n805), .B2(G322), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G179), .A2(G200), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n212), .B1(new_n807), .B2(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G294), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n212), .A2(new_n452), .A3(new_n397), .A4(G179), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n807), .A2(G20), .A3(new_n452), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n328), .B1(new_n816), .B2(G329), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n212), .A2(new_n397), .A3(G179), .A4(G190), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n817), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n798), .A2(G200), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n452), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n814), .B(new_n821), .C1(G326), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(G190), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT33), .B(G317), .Z(new_n827));
  OAI211_X1 g0627(.A(new_n806), .B(new_n824), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G58), .A2(new_n805), .B1(new_n803), .B2(new_n376), .ZN(new_n829));
  INV_X1    g0629(.A(G159), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n815), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT32), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n812), .A2(new_n470), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n820), .A2(new_n545), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n808), .A2(new_n486), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n833), .A2(new_n834), .A3(new_n255), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G50), .A2(new_n823), .B1(new_n825), .B2(G68), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n829), .A2(new_n832), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n797), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n796), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n792), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n703), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n778), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  NOR2_X1   g0644(.A1(new_n395), .A2(new_n698), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n398), .B1(new_n384), .B2(new_n719), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n395), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n691), .B2(new_n698), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n399), .A2(new_n719), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n668), .B2(new_n689), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n770), .A2(G330), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n776), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n805), .A2(G143), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G137), .A2(new_n823), .B1(new_n825), .B2(G150), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n859), .B(new_n860), .C1(new_n830), .C2(new_n802), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT100), .Z(new_n862));
  AND2_X1   g0662(.A1(new_n862), .A2(KEYINPUT34), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n811), .A2(G50), .B1(new_n819), .B2(G68), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT101), .Z(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n328), .B1(new_n815), .B2(new_n866), .C1(new_n201), .C2(new_n808), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(KEYINPUT34), .B2(new_n862), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n328), .B(new_n835), .C1(G311), .C2(new_n816), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n870), .B1(new_n470), .B2(new_n820), .C1(new_n545), .C2(new_n812), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G303), .B2(new_n823), .ZN(new_n872));
  AOI22_X1  g0672(.A1(G116), .A2(new_n803), .B1(new_n805), .B2(G294), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(new_n818), .C2(new_n826), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n797), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n790), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n797), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n849), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n779), .B1(G77), .B2(new_n877), .C1(new_n878), .C2(new_n791), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n857), .A2(new_n858), .B1(new_n875), .B2(new_n879), .ZN(G384));
  OR2_X1    g0680(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(G116), .A3(new_n220), .A4(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT36), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n376), .A2(G50), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n885), .A2(new_n408), .B1(G50), .B2(new_n202), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(G1), .A3(new_n314), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT102), .Z(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n696), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n421), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n442), .A2(new_n892), .A3(new_n893), .A4(new_n456), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n456), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n421), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n900), .B2(new_n441), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT104), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT104), .B1(new_n418), .B2(new_n420), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n891), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(new_n906), .A3(new_n891), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n895), .B1(new_n908), .B2(KEYINPUT37), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n649), .B1(KEYINPUT79), .B2(new_n460), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n910), .A2(new_n447), .B1(new_n907), .B2(new_n905), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n890), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n894), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n905), .A2(new_n907), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n890), .B1(new_n462), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n767), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT31), .B1(new_n762), .B2(new_n698), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n849), .B1(new_n921), .B2(new_n748), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n320), .A2(new_n698), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n321), .A2(new_n324), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n324), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n320), .B(new_n698), .C1(new_n296), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n889), .B1(new_n918), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n458), .B(new_n455), .C1(new_n650), .C2(new_n460), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n451), .A2(new_n696), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n252), .B1(new_n434), .B2(new_n438), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n429), .B2(new_n428), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n456), .B1(new_n451), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n935), .B2(new_n931), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n894), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT106), .B1(new_n938), .B2(new_n890), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT106), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n940), .B(KEYINPUT38), .C1(new_n932), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n462), .A2(new_n915), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT38), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n939), .A2(new_n941), .B1(new_n909), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n944), .A2(KEYINPUT40), .A3(new_n927), .A4(new_n922), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n929), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n921), .A2(new_n748), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n463), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n705), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT103), .ZN(new_n951));
  INV_X1    g0751(.A(new_n851), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n845), .B1(new_n690), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n924), .A2(new_n926), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n927), .B(KEYINPUT103), .C1(new_n852), .C2(new_n845), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n912), .A2(new_n917), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n444), .A2(new_n446), .A3(new_n696), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n912), .A2(new_n917), .A3(KEYINPUT39), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n296), .A2(new_n320), .A3(new_n719), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n931), .A2(new_n930), .B1(new_n936), .B2(new_n894), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n940), .B1(new_n963), .B2(KEYINPUT38), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n938), .A2(KEYINPUT106), .A3(new_n890), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n964), .A2(new_n965), .B1(new_n914), .B2(new_n916), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n960), .B(new_n962), .C1(KEYINPUT39), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n958), .A2(new_n959), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n463), .B1(new_n746), .B2(new_n745), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n652), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n950), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n211), .B2(new_n773), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n950), .A2(new_n971), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n884), .B(new_n888), .C1(new_n973), .C2(new_n974), .ZN(G367));
  NAND2_X1  g0775(.A1(new_n736), .A2(new_n739), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n719), .B1(new_n553), .B2(new_n564), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n976), .A2(new_n977), .B1(new_n677), .B2(new_n719), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n687), .B1(new_n978), .B2(new_n715), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(new_n698), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n677), .A2(new_n719), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n736), .A2(new_n739), .ZN(new_n982));
  INV_X1    g0782(.A(new_n977), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n615), .A2(new_n617), .A3(new_n701), .A4(new_n719), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT42), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n984), .A2(KEYINPUT42), .A3(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n980), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n490), .A2(new_n698), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n674), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n654), .B2(new_n989), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT107), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n988), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n987), .A2(new_n986), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n997), .A2(new_n993), .A3(new_n980), .A4(new_n992), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n709), .A2(new_n717), .A3(new_n978), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n996), .B2(new_n998), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n725), .B(KEYINPUT41), .Z(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n722), .B2(new_n978), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n985), .B1(new_n610), .B2(new_n698), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n984), .A2(new_n1007), .A3(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n984), .B2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n718), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n714), .A2(new_n716), .A3(new_n720), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n985), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n709), .B(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1009), .A2(new_n718), .A3(new_n1013), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1015), .A2(new_n771), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1004), .B1(new_n1020), .B2(new_n771), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1003), .B1(new_n1021), .B2(new_n775), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n992), .A2(new_n792), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n812), .A2(new_n201), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n255), .B(new_n1024), .C1(G137), .C2(new_n816), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n825), .A2(G159), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n823), .A2(G143), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n808), .A2(new_n202), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n376), .B2(new_n819), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G150), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n207), .A2(new_n802), .B1(new_n804), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n255), .B1(new_n815), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n820), .A2(new_n486), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G107), .C2(new_n809), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G294), .A2(new_n825), .B1(new_n823), .B2(G311), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n812), .B2(new_n629), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n818), .A2(new_n802), .B1(new_n804), .B2(new_n813), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1030), .A2(new_n1032), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n797), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n784), .A2(new_n242), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(new_n794), .C1(new_n215), .C2(new_n378), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n779), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT108), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1023), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1022), .A2(new_n1051), .ZN(G387));
  AOI22_X1  g0852(.A1(G311), .A2(new_n825), .B1(new_n823), .B2(G322), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n813), .B2(new_n802), .C1(new_n1033), .C2(new_n804), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n811), .A2(G294), .B1(new_n809), .B2(G283), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT110), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n820), .A2(new_n629), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n328), .B(new_n1064), .C1(G326), .C2(new_n816), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n352), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n803), .A2(G68), .B1(new_n1067), .B2(new_n825), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT109), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n255), .B(new_n1035), .C1(G150), .C2(new_n816), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n376), .A2(new_n811), .B1(new_n809), .B2(new_n379), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n823), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1071), .C1(new_n830), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n805), .B2(G50), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n797), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n717), .A2(new_n841), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n727), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n780), .A2(new_n1078), .B1(new_n545), .B2(new_n724), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n348), .A2(G50), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT50), .ZN(new_n1081));
  AOI21_X1  g0881(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n727), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n784), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n239), .A2(new_n786), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n794), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n779), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1076), .A2(new_n1077), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n775), .B2(new_n1018), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n771), .A2(new_n1018), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n725), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n771), .A2(new_n1018), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(G393));
  NOR2_X1   g0894(.A1(new_n1015), .A2(KEYINPUT111), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT111), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1019), .B1(new_n1014), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n984), .A2(new_n792), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n794), .B1(new_n486), .B2(new_n215), .C1(new_n785), .C2(new_n250), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n779), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n805), .A2(G311), .B1(G317), .B2(new_n823), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  AOI211_X1 g0903(.A(new_n328), .B(new_n834), .C1(G322), .C2(new_n816), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n811), .A2(G283), .B1(new_n809), .B2(G116), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n813), .C2(new_n826), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n803), .B2(G294), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1031), .A2(new_n1072), .B1(new_n804), .B2(new_n830), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n820), .A2(new_n470), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n255), .B(new_n1112), .C1(G143), .C2(new_n816), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n811), .A2(G68), .B1(new_n809), .B2(G77), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n207), .C2(new_n826), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n803), .B2(new_n381), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1108), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1101), .B1(new_n1119), .B2(new_n793), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1098), .A2(new_n775), .B1(new_n1099), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1091), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n725), .A3(new_n1020), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(G390));
  NAND3_X1  g0924(.A1(new_n922), .A2(new_n927), .A3(G330), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT39), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n944), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n927), .B1(new_n852), .B2(new_n845), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1128), .A2(new_n960), .B1(new_n1129), .B2(new_n961), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n744), .A2(new_n719), .A3(new_n848), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n846), .B1(new_n924), .B2(new_n926), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1132), .A2(new_n962), .A3(new_n966), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1126), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n961), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n960), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n964), .A2(new_n965), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT39), .B1(new_n1137), .B2(new_n917), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(new_n846), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n961), .B(new_n944), .C1(new_n1141), .C2(new_n954), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n927), .A2(new_n770), .A3(G330), .A4(new_n878), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1134), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n463), .A2(G330), .A3(new_n947), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n969), .A2(new_n652), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n769), .A2(new_n763), .A3(new_n766), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n741), .A2(new_n667), .A3(new_n719), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n645), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n878), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n954), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1125), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n953), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n922), .A2(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n954), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1147), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1145), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1134), .A2(new_n1159), .A3(new_n1144), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n725), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1134), .A2(new_n775), .A3(new_n1144), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n779), .B1(new_n1067), .B2(new_n877), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n328), .B(new_n833), .C1(G294), .C2(new_n816), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n809), .A2(G77), .B1(new_n819), .B2(G68), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n545), .B2(new_n826), .C1(new_n818), .C2(new_n1072), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n486), .A2(new_n802), .B1(new_n804), .B2(new_n629), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n255), .B1(new_n816), .B2(G125), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n830), .B2(new_n808), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G50), .B2(new_n819), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n811), .A2(G150), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT53), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n823), .A2(G128), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n825), .A2(G137), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT54), .B(G143), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n866), .A2(new_n804), .B1(new_n802), .B2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1169), .A2(new_n1170), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1165), .B1(new_n1181), .B2(new_n793), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1128), .A2(new_n960), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1184), .B2(new_n791), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1163), .A2(new_n1164), .A3(new_n1185), .ZN(G378));
  AOI21_X1  g0986(.A(new_n889), .B1(new_n1137), .B2(new_n917), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n922), .A2(new_n927), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n705), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n361), .A2(new_n370), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n364), .A2(new_n891), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1189), .A2(new_n929), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1189), .B2(new_n929), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n968), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n958), .A2(new_n959), .A3(new_n967), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1192), .B(new_n1193), .Z(new_n1199));
  NAND2_X1  g0999(.A1(new_n945), .A2(G330), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT40), .B1(new_n1188), .B2(new_n957), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1189), .A2(new_n929), .A3(new_n1194), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1197), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1147), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1162), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1207), .A3(KEYINPUT57), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n725), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT116), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1205), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1197), .A2(new_n1204), .A3(KEYINPUT116), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1209), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n775), .A3(new_n1213), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1194), .A2(new_n791), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n776), .B1(G50), .B2(new_n877), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n328), .A2(G41), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1028), .B(new_n1219), .C1(G283), .C2(new_n816), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n811), .A2(new_n376), .B1(new_n819), .B2(G58), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n486), .B2(new_n826), .C1(new_n629), .C2(new_n1072), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n545), .A2(new_n804), .B1(new_n802), .B2(new_n378), .ZN(new_n1224));
  XOR2_X1   g1024(.A(KEYINPUT113), .B(KEYINPUT58), .Z(new_n1225));
  OR3_X1    g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1219), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n816), .C2(G124), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n823), .A2(G125), .B1(G150), .B2(new_n809), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n866), .B2(new_n826), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1179), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n811), .A2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT114), .Z(new_n1235));
  INV_X1    g1035(.A(G128), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n804), .B2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT115), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1232), .B(new_n1238), .C1(G137), .C2(new_n803), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT59), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1230), .B1(new_n830), .B2(new_n820), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1229), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1218), .B1(new_n1244), .B2(new_n793), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1217), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1216), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT117), .B1(new_n1215), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT117), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1246), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1197), .A2(new_n1204), .A3(KEYINPUT116), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT116), .B1(new_n1197), .B2(new_n1204), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1250), .B1(new_n1253), .B2(new_n775), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1207), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1249), .B(new_n1254), .C1(new_n1255), .C2(new_n1209), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1248), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G375));
  NAND2_X1  g1058(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n775), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n779), .B1(G68), .B2(new_n877), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT118), .ZN(new_n1262));
  INV_X1    g1062(.A(G77), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n255), .B1(new_n820), .B2(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n826), .A2(new_n629), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n803), .A2(G107), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n805), .A2(G283), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n809), .A2(new_n379), .B1(new_n816), .B2(G303), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n486), .B2(new_n812), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(G294), .B2(new_n823), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G137), .A2(new_n805), .B1(new_n803), .B2(G150), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n812), .A2(new_n830), .B1(new_n207), .B2(new_n808), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n328), .B1(new_n1236), .B2(new_n815), .C1(new_n820), .C2(new_n201), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(new_n825), .C2(new_n1233), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1273), .B(new_n1276), .C1(new_n866), .C2(new_n1072), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1272), .A2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1278), .A2(KEYINPUT119), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n797), .B1(new_n1278), .B2(KEYINPUT119), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1261), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n927), .B2(new_n876), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1260), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT120), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT120), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1260), .A2(new_n1285), .A3(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1004), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1155), .A2(new_n1147), .A3(new_n1158), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1160), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(G381));
  INV_X1    g1092(.A(KEYINPUT121), .ZN(new_n1293));
  AND4_X1   g1093(.A1(new_n1022), .A2(new_n1051), .A3(new_n1123), .A4(new_n1121), .ZN(new_n1294));
  INV_X1    g1094(.A(G378), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1090), .B(new_n843), .C1(new_n1093), .C2(new_n1092), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(G384), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1294), .A2(new_n1295), .A3(new_n1291), .A4(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1293), .B1(new_n1257), .B2(new_n1299), .ZN(new_n1300));
  AOI211_X1 g1100(.A(KEYINPUT121), .B(new_n1298), .C1(new_n1248), .C2(new_n1256), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(G407));
  NAND2_X1  g1103(.A1(new_n1214), .A2(new_n1210), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1209), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1249), .B1(new_n1306), .B2(new_n1254), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1215), .A2(KEYINPUT117), .A3(new_n1247), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1295), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G213), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(G343), .ZN(new_n1311));
  XOR2_X1   g1111(.A(new_n1311), .B(KEYINPUT122), .Z(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(G213), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT123), .B1(new_n1302), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G378), .B1(new_n1248), .B2(new_n1256), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1310), .B1(new_n1316), .B2(new_n1312), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT123), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1317), .B(new_n1318), .C1(new_n1301), .C2(new_n1300), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1315), .A2(new_n1319), .ZN(G409));
  INV_X1    g1120(.A(new_n1311), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1215), .A2(new_n1295), .A3(new_n1247), .ZN(new_n1322));
  OR2_X1    g1122(.A1(new_n1205), .A2(KEYINPUT124), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n774), .B1(new_n1205), .B2(KEYINPUT124), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1250), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1212), .A2(new_n1288), .A3(new_n1207), .A4(new_n1213), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G378), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1321), .B1(new_n1322), .B2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1159), .A2(new_n726), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1155), .A2(new_n1158), .A3(new_n1147), .A4(KEYINPUT60), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT60), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1289), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1329), .A2(new_n1330), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1329), .A2(KEYINPUT125), .A3(new_n1330), .A4(new_n1332), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1287), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(G384), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1287), .A2(new_n1335), .A3(G384), .A4(new_n1336), .ZN(new_n1340));
  AOI22_X1  g1140(.A1(new_n1339), .A2(new_n1340), .B1(G2897), .B2(new_n1312), .ZN(new_n1341));
  AND4_X1   g1141(.A1(G2897), .A2(new_n1339), .A3(new_n1311), .A4(new_n1340), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1328), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1321), .B(new_n1345), .C1(new_n1322), .C2(new_n1327), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1306), .A2(G378), .A3(new_n1254), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1295), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1312), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1352), .A2(KEYINPUT63), .A3(new_n1345), .ZN(new_n1353));
  OR2_X1    g1153(.A1(G387), .A2(G390), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G393), .A2(G396), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1296), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G387), .A2(G390), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1354), .A2(new_n1356), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1356), .B1(new_n1354), .B2(new_n1357), .ZN(new_n1359));
  NOR3_X1   g1159(.A1(new_n1358), .A2(new_n1359), .A3(KEYINPUT61), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1343), .A2(new_n1348), .A3(new_n1353), .A4(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT61), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1342), .A2(new_n1341), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1362), .B1(new_n1352), .B2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1346), .A2(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1352), .A2(KEYINPUT62), .A3(new_n1345), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1364), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT126), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1369), .B(new_n1370), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1361), .B1(new_n1368), .B2(new_n1371), .ZN(G405));
  AOI21_X1  g1172(.A(new_n1295), .B1(new_n1306), .B2(new_n1254), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1309), .A2(new_n1344), .A3(new_n1374), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1345), .B1(new_n1316), .B2(new_n1373), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1375), .A2(new_n1369), .A3(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1369), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1377), .A2(new_n1378), .ZN(G402));
endmodule


