

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  XNOR2_X1 U322 ( .A(n426), .B(KEYINPUT116), .ZN(n427) );
  XNOR2_X1 U323 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U324 ( .A(n441), .B(n391), .ZN(n392) );
  XNOR2_X1 U325 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n436) );
  XOR2_X1 U326 ( .A(n404), .B(n431), .Z(n547) );
  XOR2_X1 U327 ( .A(n448), .B(n447), .Z(n516) );
  XNOR2_X1 U328 ( .A(n403), .B(n402), .ZN(n431) );
  XNOR2_X1 U329 ( .A(n428), .B(n427), .ZN(n435) );
  XNOR2_X1 U330 ( .A(n437), .B(n436), .ZN(n526) );
  XNOR2_X1 U331 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U332 ( .A(KEYINPUT28), .B(n463), .Z(n520) );
  XOR2_X1 U333 ( .A(n309), .B(n308), .Z(n563) );
  XNOR2_X1 U334 ( .A(n454), .B(G176GAT), .ZN(n455) );
  XNOR2_X1 U335 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n291) );
  XNOR2_X1 U337 ( .A(G43GAT), .B(G190GAT), .ZN(n290) );
  XNOR2_X1 U338 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U339 ( .A(n292), .B(G99GAT), .Z(n294) );
  XOR2_X1 U340 ( .A(G120GAT), .B(G71GAT), .Z(n397) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(n397), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n300) );
  XOR2_X1 U343 ( .A(G183GAT), .B(KEYINPUT19), .Z(n296) );
  XNOR2_X1 U344 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n448) );
  XOR2_X1 U346 ( .A(G15GAT), .B(n448), .Z(n298) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U349 ( .A(n300), .B(n299), .Z(n309) );
  XNOR2_X1 U350 ( .A(G127GAT), .B(KEYINPUT83), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n301), .B(KEYINPUT0), .ZN(n302) );
  XOR2_X1 U352 ( .A(n302), .B(KEYINPUT84), .Z(n304) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(G134GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n327) );
  XOR2_X1 U355 ( .A(G176GAT), .B(KEYINPUT87), .Z(n306) );
  XNOR2_X1 U356 ( .A(KEYINPUT85), .B(KEYINPUT67), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n327), .B(n307), .ZN(n308) );
  INV_X1 U359 ( .A(n563), .ZN(n453) );
  XOR2_X1 U360 ( .A(G57GAT), .B(G155GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(G1GAT), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U363 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT95), .B(KEYINPUT6), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U367 ( .A(KEYINPUT4), .B(KEYINPUT96), .Z(n317) );
  NAND2_X1 U368 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U370 ( .A(KEYINPUT94), .B(n318), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U372 ( .A(G85GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(G162GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U376 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n326) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n339) );
  XNOR2_X1 U379 ( .A(n327), .B(n339), .ZN(n328) );
  XOR2_X1 U380 ( .A(n329), .B(n328), .Z(n569) );
  XNOR2_X1 U381 ( .A(G78GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n330), .B(G148GAT), .ZN(n396) );
  XOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .Z(n410) );
  XOR2_X1 U384 ( .A(n396), .B(n410), .Z(n332) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n343) );
  XOR2_X1 U387 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n334) );
  XNOR2_X1 U388 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n335), .B(G106GAT), .Z(n337) );
  XOR2_X1 U391 ( .A(G22GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U392 ( .A(n357), .B(G218GAT), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U394 ( .A(n338), .B(KEYINPUT23), .Z(n341) );
  XNOR2_X1 U395 ( .A(n339), .B(KEYINPUT24), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U398 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n345) );
  XNOR2_X1 U399 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U401 ( .A(G197GAT), .B(n346), .ZN(n443) );
  XNOR2_X1 U402 ( .A(n347), .B(n443), .ZN(n463) );
  AND2_X1 U403 ( .A1(n569), .A2(n463), .ZN(n451) );
  XOR2_X1 U404 ( .A(KEYINPUT79), .B(KEYINPUT82), .Z(n349) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U407 ( .A(KEYINPUT15), .B(G64GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U410 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U411 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n355) );
  XNOR2_X1 U412 ( .A(G183GAT), .B(KEYINPUT80), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U416 ( .A(G78GAT), .B(G211GAT), .Z(n361) );
  XNOR2_X1 U417 ( .A(G127GAT), .B(G71GAT), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U419 ( .A(n363), .B(n362), .Z(n365) );
  XOR2_X1 U420 ( .A(G15GAT), .B(G1GAT), .Z(n380) );
  XOR2_X1 U421 ( .A(G57GAT), .B(KEYINPUT13), .Z(n395) );
  XNOR2_X1 U422 ( .A(n380), .B(n395), .ZN(n364) );
  XOR2_X1 U423 ( .A(n365), .B(n364), .Z(n581) );
  INV_X1 U424 ( .A(n581), .ZN(n557) );
  XOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n367) );
  NAND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U428 ( .A(n368), .B(KEYINPUT68), .Z(n376) );
  XOR2_X1 U429 ( .A(G22GAT), .B(G141GAT), .Z(n370) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(G36GAT), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U432 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n372) );
  XNOR2_X1 U433 ( .A(G197GAT), .B(G113GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U437 ( .A(G169GAT), .B(G8GAT), .Z(n444) );
  XOR2_X1 U438 ( .A(n377), .B(n444), .Z(n382) );
  XOR2_X1 U439 ( .A(G29GAT), .B(G43GAT), .Z(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n420) );
  XNOR2_X1 U442 ( .A(n420), .B(n380), .ZN(n381) );
  XOR2_X1 U443 ( .A(n382), .B(n381), .Z(n573) );
  INV_X1 U444 ( .A(n573), .ZN(n555) );
  XNOR2_X1 U445 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n404) );
  XOR2_X1 U446 ( .A(KEYINPUT71), .B(G85GAT), .Z(n384) );
  XNOR2_X1 U447 ( .A(G99GAT), .B(G106GAT), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n411) );
  XNOR2_X1 U449 ( .A(n411), .B(KEYINPUT32), .ZN(n388) );
  INV_X1 U450 ( .A(n388), .ZN(n386) );
  AND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  INV_X1 U452 ( .A(n387), .ZN(n385) );
  NAND2_X1 U453 ( .A1(n386), .A2(n385), .ZN(n390) );
  NAND2_X1 U454 ( .A1(n388), .A2(n387), .ZN(n389) );
  NAND2_X1 U455 ( .A1(n390), .A2(n389), .ZN(n393) );
  XOR2_X1 U456 ( .A(G176GAT), .B(G64GAT), .Z(n441) );
  XOR2_X1 U457 ( .A(G92GAT), .B(KEYINPUT73), .Z(n391) );
  XOR2_X1 U458 ( .A(n395), .B(n394), .Z(n403) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U460 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n399) );
  XNOR2_X1 U461 ( .A(KEYINPUT74), .B(KEYINPUT72), .ZN(n398) );
  XOR2_X1 U462 ( .A(n399), .B(n398), .Z(n400) );
  NAND2_X1 U463 ( .A1(n555), .A2(n547), .ZN(n405) );
  XOR2_X1 U464 ( .A(n405), .B(KEYINPUT46), .Z(n406) );
  NOR2_X1 U465 ( .A1(n557), .A2(n406), .ZN(n407) );
  XNOR2_X1 U466 ( .A(KEYINPUT114), .B(n407), .ZN(n425) );
  XOR2_X1 U467 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n409) );
  XNOR2_X1 U468 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n424) );
  XOR2_X1 U470 ( .A(n411), .B(n410), .Z(n413) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U473 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n415) );
  XNOR2_X1 U474 ( .A(KEYINPUT75), .B(KEYINPUT77), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U477 ( .A(G92GAT), .B(G218GAT), .Z(n419) );
  XNOR2_X1 U478 ( .A(G36GAT), .B(G190GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n438) );
  XNOR2_X1 U480 ( .A(n420), .B(n438), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n553) );
  NAND2_X1 U483 ( .A1(n425), .A2(n553), .ZN(n428) );
  XOR2_X1 U484 ( .A(KEYINPUT47), .B(KEYINPUT115), .Z(n426) );
  XOR2_X1 U485 ( .A(KEYINPUT78), .B(n553), .Z(n562) );
  XOR2_X1 U486 ( .A(KEYINPUT36), .B(n562), .Z(n584) );
  NOR2_X1 U487 ( .A1(n584), .A2(n581), .ZN(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT45), .B(KEYINPUT117), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n433) );
  BUF_X1 U490 ( .A(n431), .Z(n578) );
  NAND2_X1 U491 ( .A1(n578), .A2(n573), .ZN(n432) );
  NOR2_X1 U492 ( .A1(n433), .A2(n432), .ZN(n434) );
  NOR2_X1 U493 ( .A1(n435), .A2(n434), .ZN(n437) );
  XOR2_X1 U494 ( .A(n438), .B(G204GAT), .Z(n440) );
  NAND2_X1 U495 ( .A1(G226GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U497 ( .A(n442), .B(n441), .Z(n446) );
  XOR2_X1 U498 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  INV_X1 U500 ( .A(n516), .ZN(n449) );
  NOR2_X1 U501 ( .A1(n526), .A2(n449), .ZN(n450) );
  XNOR2_X1 U502 ( .A(KEYINPUT54), .B(n450), .ZN(n568) );
  AND2_X1 U503 ( .A1(n451), .A2(n568), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n452), .B(KEYINPUT55), .ZN(n565) );
  NOR2_X1 U505 ( .A1(n453), .A2(n565), .ZN(n558) );
  NAND2_X1 U506 ( .A1(n558), .A2(n547), .ZN(n456) );
  XOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n474) );
  NAND2_X1 U509 ( .A1(n555), .A2(n578), .ZN(n488) );
  NOR2_X1 U510 ( .A1(n562), .A2(n581), .ZN(n457) );
  XNOR2_X1 U511 ( .A(KEYINPUT16), .B(n457), .ZN(n472) );
  INV_X1 U512 ( .A(n520), .ZN(n530) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(KEYINPUT97), .Z(n458) );
  XOR2_X1 U514 ( .A(n516), .B(n458), .Z(n525) );
  NOR2_X1 U515 ( .A1(n525), .A2(n563), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n530), .A2(n459), .ZN(n460) );
  INV_X1 U517 ( .A(n569), .ZN(n528) );
  NAND2_X1 U518 ( .A1(n460), .A2(n528), .ZN(n470) );
  NAND2_X1 U519 ( .A1(n516), .A2(n563), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n463), .A2(n461), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n462), .Z(n466) );
  NOR2_X1 U522 ( .A1(n463), .A2(n563), .ZN(n464) );
  XOR2_X1 U523 ( .A(n464), .B(KEYINPUT26), .Z(n570) );
  OR2_X1 U524 ( .A1(n570), .A2(n525), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U526 ( .A(KEYINPUT98), .B(n467), .Z(n468) );
  NAND2_X1 U527 ( .A1(n468), .A2(n569), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n484) );
  INV_X1 U529 ( .A(n484), .ZN(n471) );
  NAND2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n503) );
  NOR2_X1 U531 ( .A1(n488), .A2(n503), .ZN(n479) );
  NAND2_X1 U532 ( .A1(n479), .A2(n528), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n479), .A2(n516), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U538 ( .A1(n479), .A2(n563), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n520), .A2(n479), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT100), .ZN(n481) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n483) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n492) );
  NOR2_X1 U546 ( .A1(n557), .A2(n484), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n485), .B(KEYINPUT101), .ZN(n486) );
  NOR2_X1 U548 ( .A1(n584), .A2(n486), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n487), .ZN(n514) );
  NOR2_X1 U550 ( .A1(n514), .A2(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n500) );
  NAND2_X1 U553 ( .A1(n500), .A2(n528), .ZN(n491) );
  XOR2_X1 U554 ( .A(n492), .B(n491), .Z(G1328GAT) );
  XOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT105), .Z(n494) );
  NAND2_X1 U556 ( .A1(n500), .A2(n516), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n496) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(KEYINPUT107), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n563), .A2(n500), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n497), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n500), .A2(n520), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  NAND2_X1 U567 ( .A1(n547), .A2(n573), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT109), .B(n502), .Z(n513) );
  NOR2_X1 U569 ( .A1(n513), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(KEYINPUT110), .B(n504), .ZN(n510) );
  NAND2_X1 U571 ( .A1(n528), .A2(n510), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n516), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT111), .Z(n509) );
  NAND2_X1 U576 ( .A1(n510), .A2(n563), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U579 ( .A1(n510), .A2(n520), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n528), .A2(n521), .ZN(n515) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n563), .A2(n521), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n518), .B(KEYINPUT112), .ZN(n519) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n523) );
  NAND2_X1 U590 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT119), .Z(n533) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(KEYINPUT118), .B(n529), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n530), .A2(n563), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n541), .A2(n531), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n538), .A2(n555), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U602 ( .A1(n538), .A2(n547), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n557), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U608 ( .A1(n538), .A2(n562), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT120), .ZN(n543) );
  NOR2_X1 U611 ( .A1(n570), .A2(n541), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n555), .A2(n551), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n545) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n544) );
  XNOR2_X1 U616 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U617 ( .A(KEYINPUT52), .B(n546), .Z(n549) );
  NAND2_X1 U618 ( .A1(n551), .A2(n547), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n551), .A2(n557), .ZN(n550) );
  XNOR2_X1 U621 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U622 ( .A(n551), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U625 ( .A1(n555), .A2(n558), .ZN(n556) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  OR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  AND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n572) );
  INV_X1 U636 ( .A(n570), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n583) );
  NOR2_X1 U638 ( .A1(n583), .A2(n573), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G218GAT), .B(n587), .Z(G1355GAT) );
endmodule

