//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G58), .C2(G232), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G1), .B2(G20), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n219), .A2(new_n220), .A3(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n203), .A2(G50), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n218), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n208), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  INV_X1    g0041(.A(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  INV_X1    g0044(.A(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n207), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  NOR2_X1   g0049(.A1(new_n220), .A2(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G13), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G20), .A2(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT15), .B(G87), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n220), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n220), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n253), .B1(new_n254), .B2(new_n255), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n252), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n262), .A2(new_n250), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  OAI211_X1 g0072(.A(G1), .B(G13), .C1(new_n256), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(G244), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n256), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G107), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(G1698), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n282), .B(new_n286), .C1(new_n287), .C2(new_n212), .ZN(new_n288));
  INV_X1    g0088(.A(new_n273), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n271), .B(new_n276), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n267), .B1(new_n290), .B2(G169), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT73), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n292), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n280), .A2(G226), .A3(new_n281), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n289), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(G238), .A3(new_n268), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(new_n270), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT13), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n303), .A2(new_n307), .A3(new_n304), .A4(new_n270), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(KEYINPUT75), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT75), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(new_n310), .A3(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(G169), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(G179), .A3(new_n308), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n309), .A2(new_n315), .A3(G169), .A4(new_n311), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n251), .A2(KEYINPUT12), .A3(G68), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT76), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT12), .B1(new_n251), .B2(G68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G50), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n257), .A2(new_n322), .B1(new_n255), .B2(new_n264), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n220), .A2(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n262), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT11), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n262), .A2(new_n250), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n321), .B(new_n326), .C1(new_n211), .C2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n298), .B1(new_n317), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G226), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n270), .B1(new_n274), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n332), .A2(KEYINPUT68), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n264), .B2(new_n280), .ZN(new_n336));
  INV_X1    g0136(.A(new_n287), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(G223), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n333), .B(new_n334), .C1(new_n338), .C2(new_n273), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(KEYINPUT69), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G190), .ZN(new_n343));
  OAI21_X1  g0143(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n344));
  INV_X1    g0144(.A(G150), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT8), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n242), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT70), .B(G58), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n344), .B1(new_n345), .B2(new_n257), .C1(new_n349), .C2(new_n255), .ZN(new_n350));
  INV_X1    g0150(.A(new_n251), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n262), .B1(new_n322), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n322), .B2(new_n328), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(KEYINPUT74), .B2(KEYINPUT9), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n340), .A2(G200), .A3(new_n341), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n343), .A2(new_n357), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT10), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n356), .B(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT10), .A3(new_n343), .A4(new_n358), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n340), .A2(new_n341), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n353), .C1(G179), .C2(new_n366), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n309), .A2(G200), .A3(new_n311), .ZN(new_n371));
  INV_X1    g0171(.A(new_n329), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n306), .A2(G190), .A3(new_n308), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n252), .B(new_n265), .C1(new_n259), .C2(new_n262), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT71), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n290), .A2(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT72), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n290), .A2(G190), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n288), .A2(new_n289), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n270), .ZN(new_n385));
  OAI21_X1  g0185(.A(G200), .B1(new_n385), .B2(new_n276), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n378), .A2(new_n379), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT72), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n256), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT77), .A2(G33), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(KEYINPUT3), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n278), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT7), .B1(new_n396), .B2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n395), .A2(new_n398), .A3(new_n220), .A4(new_n278), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G68), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G159), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n257), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(KEYINPUT70), .A2(G58), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT70), .A2(G58), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n202), .B1(new_n405), .B2(G68), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n407), .B2(G20), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AND2_X1   g0210(.A1(KEYINPUT77), .A2(G33), .ZN(new_n411));
  NOR2_X1   g0211(.A1(KEYINPUT77), .A2(G33), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n277), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n413), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n279), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n398), .B1(new_n280), .B2(G20), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n211), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n406), .A2(new_n220), .B1(new_n401), .B2(new_n257), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n410), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(new_n262), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n328), .A2(new_n349), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n351), .B2(new_n349), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n273), .A2(G232), .A3(new_n268), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n270), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n270), .A3(KEYINPUT78), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n281), .A2(G226), .ZN(new_n428));
  NOR2_X1   g0228(.A1(G223), .A2(G1698), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n428), .B(new_n429), .C1(new_n395), .C2(new_n278), .ZN(new_n430));
  INV_X1    g0230(.A(G87), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n256), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n289), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G200), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n433), .A3(G190), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n419), .A2(new_n421), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n419), .A2(new_n421), .ZN(new_n440));
  INV_X1    g0240(.A(new_n428), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n396), .B(new_n441), .C1(G223), .C2(G1698), .ZN(new_n442));
  INV_X1    g0242(.A(new_n432), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n273), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n422), .A2(KEYINPUT78), .A3(new_n270), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT78), .B1(new_n422), .B2(new_n270), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G169), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n294), .B2(new_n434), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT18), .B1(new_n440), .B2(new_n449), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n438), .A2(new_n439), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AND4_X1   g0253(.A1(new_n330), .A2(new_n376), .A3(new_n391), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n262), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n219), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n251), .A3(G116), .A4(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n260), .A2(new_n261), .B1(G20), .B2(new_n207), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n220), .C1(G33), .C2(new_n213), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n458), .A2(KEYINPUT20), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT20), .B1(new_n458), .B2(new_n460), .ZN(new_n462));
  OAI221_X1 g0262(.A(new_n457), .B1(G116), .B2(new_n251), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G179), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n273), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n208), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n466), .B(G274), .C1(new_n468), .C2(new_n467), .ZN(new_n473));
  INV_X1    g0273(.A(G303), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n280), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G257), .A2(G1698), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n395), .B2(new_n278), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n281), .A2(G264), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n472), .B(new_n473), .C1(new_n479), .C2(new_n273), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n464), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n463), .A2(G169), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT21), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n480), .A2(new_n485), .A3(G169), .A4(new_n463), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n481), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n463), .B1(new_n480), .B2(G200), .ZN(new_n488));
  INV_X1    g0288(.A(new_n479), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n289), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n490), .A2(G190), .A3(new_n472), .A4(new_n473), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT85), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT85), .B1(new_n488), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n487), .B(new_n496), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n431), .A2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n396), .A2(KEYINPUT22), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n411), .A2(new_n412), .A3(new_n207), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n283), .B2(new_n284), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n220), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n220), .A2(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT23), .ZN(new_n507));
  NAND2_X1  g0307(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n508));
  NOR2_X1   g0308(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n500), .A2(new_n504), .A3(new_n507), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n509), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n262), .A3(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n455), .A2(new_n251), .A3(new_n456), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n251), .A2(G107), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT25), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n469), .A2(G264), .A3(new_n273), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n411), .A2(new_n412), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n395), .B2(new_n278), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n281), .A2(G257), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n473), .B(new_n520), .C1(new_n527), .C2(new_n273), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G179), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n367), .B2(new_n528), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n220), .B1(new_n301), .B2(new_n533), .ZN(new_n534));
  AND4_X1   g0334(.A1(KEYINPUT82), .A2(new_n431), .A3(new_n213), .A4(new_n245), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G87), .A2(G97), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT82), .B1(new_n536), .B2(new_n245), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n533), .B1(new_n255), .B2(new_n213), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI211_X1 g0340(.A(G20), .B(new_n211), .C1(new_n395), .C2(new_n278), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n532), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n396), .A2(new_n220), .A3(G68), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(KEYINPUT83), .A3(new_n538), .A4(new_n539), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n262), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n351), .A2(new_n254), .ZN(new_n546));
  INV_X1    g0346(.A(new_n254), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n515), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n466), .A2(G274), .ZN(new_n552));
  XOR2_X1   g0352(.A(new_n552), .B(KEYINPUT81), .Z(new_n553));
  OAI211_X1 g0353(.A(new_n273), .B(G250), .C1(G1), .C2(new_n465), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n395), .A2(new_n278), .B1(new_n275), .B2(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n212), .A2(new_n281), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n501), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n553), .B(new_n554), .C1(new_n557), .C2(new_n273), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G169), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n294), .B2(new_n558), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n545), .A2(KEYINPUT84), .A3(new_n546), .A4(new_n548), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n551), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n411), .A2(new_n412), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n284), .B1(new_n563), .B2(KEYINPUT3), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n564), .A2(new_n525), .A3(new_n523), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n289), .B1(new_n565), .B2(new_n522), .ZN(new_n566));
  INV_X1    g0366(.A(G190), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n473), .A4(new_n520), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n528), .A2(new_n377), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n570), .A2(new_n514), .A3(new_n516), .A4(new_n518), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n545), .A2(new_n546), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n558), .A2(new_n567), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n515), .A2(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n558), .A2(G200), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n531), .A2(new_n562), .A3(new_n571), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n275), .A2(G1698), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n564), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n579), .B(KEYINPUT4), .C1(new_n284), .C2(new_n283), .ZN(new_n582));
  OAI211_X1 g0382(.A(G250), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(new_n459), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n273), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n473), .B1(new_n470), .B2(new_n214), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT79), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n580), .B1(new_n395), .B2(new_n278), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(KEYINPUT4), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(new_n583), .A3(new_n459), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n289), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT79), .ZN(new_n592));
  INV_X1    g0392(.A(new_n586), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G190), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n597), .A2(new_n213), .A3(G107), .ZN(new_n598));
  XNOR2_X1  g0398(.A(G97), .B(G107), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n600), .A2(new_n220), .B1(new_n264), .B2(new_n257), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n245), .B1(new_n414), .B2(new_n415), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n262), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n251), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n515), .B2(G97), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n584), .B1(KEYINPUT4), .B2(new_n588), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n586), .B1(new_n607), .B2(new_n289), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n596), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n587), .A2(new_n367), .A3(new_n594), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n608), .A2(new_n294), .B1(new_n603), .B2(new_n605), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n612), .A2(KEYINPUT80), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT80), .B1(new_n612), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n577), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n454), .A2(new_n498), .A3(new_n617), .ZN(G372));
  NAND2_X1  g0418(.A1(new_n560), .A2(new_n549), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT89), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n612), .A2(new_n613), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT80), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT80), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n624), .A2(new_n562), .A3(new_n625), .A4(new_n576), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n574), .A2(new_n575), .A3(new_n546), .A4(new_n545), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n573), .B1(new_n560), .B2(new_n549), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(new_n622), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n621), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n595), .A2(G190), .B1(G200), .B2(new_n609), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n624), .A2(new_n625), .B1(new_n606), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n576), .A2(new_n571), .A3(new_n619), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(KEYINPUT88), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n576), .A2(new_n571), .A3(new_n619), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n616), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n531), .A2(new_n487), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n454), .B1(new_n633), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n369), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n438), .A2(new_n439), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n330), .A2(new_n645), .A3(new_n375), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n450), .A2(new_n451), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n362), .A2(new_n365), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n650), .ZN(G369));
  INV_X1    g0451(.A(new_n531), .ZN(new_n652));
  INV_X1    g0452(.A(G13), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G20), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n219), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n519), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n531), .A2(new_n662), .A3(new_n571), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n495), .A2(new_n497), .B1(new_n463), .B2(new_n660), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n463), .A2(new_n660), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n487), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(G330), .B(new_n664), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n531), .A2(new_n662), .A3(new_n571), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n487), .A2(new_n660), .ZN(new_n670));
  INV_X1    g0470(.A(new_n660), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n669), .A2(new_n670), .B1(new_n652), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(G399));
  NOR2_X1   g0473(.A1(new_n535), .A2(new_n537), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n207), .ZN(new_n675));
  INV_X1    g0475(.A(new_n221), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n675), .A2(new_n219), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n680));
  INV_X1    g0480(.A(new_n677), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n679), .B(new_n680), .C1(new_n226), .C2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n683));
  XNOR2_X1  g0483(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n498), .A2(new_n617), .A3(new_n671), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n558), .A2(new_n294), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n595), .A2(new_n482), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n566), .A2(new_n520), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT30), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n482), .A2(new_n608), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n294), .A3(new_n528), .A4(new_n558), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n686), .B(new_n694), .C1(new_n688), .C2(new_n689), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n660), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n699), .A3(new_n660), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT94), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n616), .A2(new_n639), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n620), .B1(new_n705), .B2(new_n641), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n626), .A2(new_n630), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n631), .A2(new_n576), .A3(new_n619), .A4(KEYINPUT26), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n629), .A2(new_n710), .A3(KEYINPUT26), .A4(new_n631), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n704), .A2(new_n713), .A3(KEYINPUT29), .A4(new_n671), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n660), .B1(new_n706), .B2(new_n712), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n704), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n671), .B1(new_n642), .B2(new_n633), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n703), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n684), .B1(new_n721), .B2(G1), .ZN(G364));
  NOR3_X1   g0522(.A1(new_n653), .A2(new_n465), .A3(G20), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n677), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n665), .A2(new_n667), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(G330), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n728), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n280), .A2(new_n221), .A3(G355), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n243), .A2(new_n465), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n396), .A2(new_n676), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G45), .B2(new_n226), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT96), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n731), .B1(G116), .B2(new_n221), .C1(new_n732), .C2(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(KEYINPUT97), .A2(G169), .ZN(new_n737));
  NOR2_X1   g0537(.A1(KEYINPUT97), .A2(G169), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n261), .B1(new_n739), .B2(G20), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n727), .ZN(new_n746));
  NOR4_X1   g0546(.A1(new_n220), .A2(new_n294), .A3(G190), .A4(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G311), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n285), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n220), .A2(new_n294), .A3(new_n567), .A4(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n220), .B1(new_n754), .B2(G190), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n752), .A2(new_n753), .B1(new_n755), .B2(new_n521), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n294), .A2(new_n377), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G20), .A3(new_n567), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT33), .B(G317), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n750), .B(new_n756), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n220), .A2(new_n567), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n377), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G303), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT98), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n757), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(new_n757), .B2(new_n762), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G326), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT99), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n220), .B2(G190), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n567), .A2(KEYINPUT99), .A3(G20), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n763), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n774), .A2(new_n754), .A3(new_n775), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G283), .A2(new_n777), .B1(new_n779), .B2(G329), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n761), .A2(new_n766), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n755), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n405), .A2(new_n751), .B1(new_n782), .B2(G97), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n783), .B1(new_n431), .B2(new_n764), .C1(new_n770), .C2(new_n322), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n778), .A2(new_n401), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n280), .B1(new_n758), .B2(new_n211), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G77), .B2(new_n747), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(new_n245), .C2(new_n776), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n781), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n746), .B1(new_n790), .B2(new_n740), .ZN(new_n791));
  INV_X1    g0591(.A(new_n743), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n745), .B(new_n791), .C1(new_n728), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n730), .A2(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n267), .A2(new_n660), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n391), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n297), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n298), .A2(new_n795), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n718), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n799), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n671), .B(new_n801), .C1(new_n642), .C2(new_n633), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n703), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n746), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT101), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n800), .A2(new_n802), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n703), .B2(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n752), .A2(new_n521), .B1(new_n755), .B2(new_n213), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n285), .B1(new_n764), .B2(new_n245), .C1(new_n810), .C2(new_n758), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n776), .A2(new_n431), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n778), .A2(new_n749), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n809), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n814), .B1(new_n207), .B2(new_n748), .C1(new_n474), .C2(new_n770), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT100), .Z(new_n816));
  NOR2_X1   g0616(.A1(new_n764), .A2(new_n322), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n759), .A2(G150), .B1(new_n751), .B2(G143), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n401), .B2(new_n748), .C1(new_n770), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT34), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n211), .A2(new_n776), .B1(new_n778), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n564), .B(new_n825), .C1(new_n405), .C2(new_n782), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n816), .B1(new_n817), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n746), .B1(new_n828), .B2(new_n740), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n740), .A2(new_n741), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n264), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(new_n742), .C2(new_n801), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n808), .A2(new_n832), .ZN(G384));
  NAND2_X1  g0633(.A1(new_n317), .A2(new_n329), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n329), .A2(new_n660), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n374), .A3(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n329), .B(new_n660), .C1(new_n317), .C2(new_n375), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n799), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n698), .A2(new_n838), .A3(new_n700), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n409), .A2(new_n262), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n400), .A2(new_n408), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(KEYINPUT16), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n449), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n421), .A2(new_n844), .B1(new_n845), .B2(new_n658), .ZN(new_n846));
  INV_X1    g0646(.A(new_n437), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n658), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n440), .B1(new_n449), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n437), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n658), .B1(new_n844), .B2(new_n421), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n452), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n658), .B1(new_n419), .B2(new_n421), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n452), .A2(KEYINPUT103), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT103), .B1(new_n452), .B2(new_n857), .ZN(new_n859));
  INV_X1    g0659(.A(new_n852), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n851), .B1(new_n850), .B2(new_n437), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n856), .B1(new_n863), .B2(KEYINPUT38), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n698), .A2(new_n838), .A3(new_n700), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n841), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT40), .ZN(new_n870));
  INV_X1    g0670(.A(new_n856), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n853), .B2(new_n855), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n701), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n454), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G330), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n836), .A2(new_n837), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n298), .A2(new_n671), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT102), .Z(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n802), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n873), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n886), .A2(new_n887), .B1(new_n647), .B2(new_n658), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n889), .B(new_n856), .C1(new_n863), .C2(KEYINPUT38), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT39), .B1(new_n871), .B2(new_n872), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n834), .A2(new_n660), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n635), .A2(new_n641), .A3(new_n636), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n621), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT29), .B(new_n671), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT94), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n715), .A2(new_n704), .A3(KEYINPUT29), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n454), .A2(new_n720), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n650), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n895), .B(new_n903), .Z(new_n904));
  XNOR2_X1  g0704(.A(new_n880), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n219), .B2(new_n654), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT35), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n225), .B1(new_n600), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(G116), .C1(new_n907), .C2(new_n600), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n264), .B(new_n226), .C1(G68), .C2(new_n405), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n201), .A2(new_n211), .ZN(new_n912));
  OAI211_X1 g0712(.A(G1), .B(new_n653), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(new_n910), .A3(new_n913), .ZN(G367));
  INV_X1    g0714(.A(KEYINPUT108), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n606), .A2(new_n671), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n635), .A2(new_n917), .B1(new_n631), .B2(new_n660), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n668), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n669), .A2(new_n670), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT42), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT42), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n616), .A2(new_n916), .B1(new_n622), .B2(new_n671), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(new_n652), .B1(new_n624), .B2(new_n625), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n922), .B(new_n923), .C1(new_n660), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n572), .A2(new_n574), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n660), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n629), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n621), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n920), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n920), .A2(new_n926), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n935), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n937), .A2(new_n932), .B1(KEYINPUT43), .B2(new_n930), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n677), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT44), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n672), .B2(new_n924), .ZN(new_n944));
  INV_X1    g0744(.A(new_n670), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n945), .A2(new_n663), .B1(new_n531), .B2(new_n660), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n918), .A2(new_n946), .A3(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n918), .B2(new_n946), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n672), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n668), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n728), .A2(G330), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n921), .B1(new_n664), .B2(new_n670), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n728), .A2(new_n956), .A3(G330), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n948), .A2(new_n952), .A3(new_n668), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n721), .A2(new_n954), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n942), .B1(new_n962), .B2(new_n721), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n940), .B1(new_n963), .B2(new_n726), .ZN(new_n964));
  INV_X1    g0764(.A(new_n201), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n280), .B1(new_n748), .B2(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n752), .A2(new_n345), .B1(new_n755), .B2(new_n211), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(G159), .C2(new_n759), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n765), .A2(new_n405), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n771), .A2(G143), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G77), .A2(new_n777), .B1(new_n779), .B2(G137), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n748), .A2(new_n810), .B1(new_n755), .B2(new_n245), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT105), .B1(new_n764), .B2(new_n207), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(G303), .C2(new_n751), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n396), .B1(new_n779), .B2(G317), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n213), .B2(new_n776), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT106), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(KEYINPUT106), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n771), .A2(G311), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n976), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n758), .A2(new_n521), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n740), .ZN(new_n986));
  INV_X1    g0786(.A(new_n733), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n744), .B1(new_n221), .B2(new_n254), .C1(new_n237), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n727), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n792), .B2(new_n930), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n915), .B1(new_n964), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n720), .A2(new_n900), .A3(new_n901), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n877), .A2(G330), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n993), .A2(new_n960), .A3(new_n994), .A4(new_n961), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n721), .B1(new_n995), .B2(new_n953), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n726), .B1(new_n996), .B2(new_n941), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n915), .B(new_n991), .C1(new_n997), .C2(new_n939), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n992), .A2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n993), .A2(new_n994), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n960), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n993), .A2(new_n994), .A3(new_n960), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(new_n677), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n960), .A2(new_n726), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n258), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT110), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(G68), .A2(G77), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n675), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1011));
  AND4_X1   g0811(.A1(new_n465), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n234), .A2(G45), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT109), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n733), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n675), .A2(new_n221), .A3(new_n280), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n221), .A2(G107), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n744), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n751), .A2(G317), .B1(new_n747), .B2(G303), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n749), .B2(new_n758), .C1(new_n770), .C2(new_n753), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n810), .B2(new_n755), .C1(new_n521), .C2(new_n764), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n779), .A2(G326), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n396), .B1(new_n777), .B2(G116), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n349), .A2(new_n758), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G50), .A2(new_n751), .B1(new_n782), .B2(new_n547), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n211), .B2(new_n748), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G77), .B2(new_n765), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G97), .A2(new_n777), .B1(new_n779), .B2(G150), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n564), .B1(new_n771), .B2(G159), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n740), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1020), .A2(new_n1039), .A3(new_n727), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT111), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n664), .B2(new_n792), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1005), .A2(new_n1006), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1005), .A2(KEYINPUT112), .A3(new_n1006), .A4(new_n1042), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(G393));
  AOI22_X1  g0847(.A1(new_n771), .A2(G317), .B1(G311), .B2(new_n751), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT114), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n245), .A2(new_n776), .B1(new_n778), .B2(new_n753), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n285), .B1(new_n764), .B2(new_n810), .C1(new_n474), .C2(new_n758), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G116), .C2(new_n782), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1053), .C1(new_n521), .C2(new_n748), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n564), .B1(G77), .B2(new_n782), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n965), .B2(new_n758), .C1(new_n258), .C2(new_n748), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n812), .B(new_n1056), .C1(G143), .C2(new_n779), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n770), .A2(new_n345), .B1(new_n401), .B2(new_n752), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT51), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n211), .C2(new_n764), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n746), .B1(new_n1061), .B2(new_n740), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n744), .B1(new_n213), .B2(new_n221), .C1(new_n248), .C2(new_n987), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n792), .C2(new_n924), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n961), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n953), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n668), .C1(new_n948), .C2(new_n952), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n726), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n995), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1004), .A2(new_n1069), .B1(new_n1072), .B2(new_n954), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n1073), .B2(new_n677), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND4_X1  g0875(.A1(new_n698), .A2(G330), .A3(new_n700), .A4(new_n801), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1076), .A2(new_n882), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n893), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n621), .A2(new_n627), .A3(new_n632), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n660), .B(new_n799), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n881), .B1(new_n1081), .B2(new_n884), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n892), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n864), .A2(new_n1078), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n715), .A2(new_n801), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n883), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n881), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1077), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT38), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n859), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n452), .A2(KEYINPUT103), .A3(new_n857), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1089), .B1(new_n1092), .B2(new_n862), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n893), .B1(new_n1093), .B2(new_n856), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1085), .A2(new_n883), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n882), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1076), .A2(new_n882), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n886), .A2(new_n893), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(new_n892), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n454), .A2(G330), .A3(new_n877), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n902), .A2(new_n650), .A3(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1076), .A2(new_n882), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1102), .A2(new_n1077), .B1(new_n1081), .B2(new_n884), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1076), .A2(new_n882), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1097), .A2(new_n1095), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1088), .A2(new_n1099), .A3(new_n1101), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n677), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1088), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1099), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1107), .A2(KEYINPUT115), .A3(new_n677), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1110), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n830), .A2(new_n349), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n280), .B1(new_n748), .B2(new_n1119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n752), .A2(new_n824), .B1(new_n755), .B2(new_n401), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n771), .C2(G128), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n765), .A2(G150), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n965), .A2(new_n776), .B1(new_n778), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1122), .B(new_n1127), .C1(new_n819), .C2(new_n758), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n285), .B1(new_n764), .B2(new_n431), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT117), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G77), .B2(new_n782), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n752), .A2(new_n207), .B1(new_n211), .B2(new_n776), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n771), .B2(G283), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n521), .C2(new_n778), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n748), .A2(new_n213), .B1(new_n245), .B2(new_n758), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT116), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n746), .B1(new_n1137), .B2(new_n740), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1117), .B(new_n1138), .C1(new_n892), .C2(new_n742), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT118), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n726), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1116), .A2(new_n1142), .ZN(G378));
  INV_X1    g0943(.A(KEYINPUT56), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n353), .A2(new_n849), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n370), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT55), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n362), .A2(new_n365), .A3(new_n369), .A4(new_n1145), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT55), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT56), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n741), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n830), .A2(new_n965), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n770), .A2(new_n1125), .B1(new_n345), .B2(new_n755), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT120), .Z(new_n1161));
  OAI22_X1  g0961(.A1(new_n748), .A2(new_n819), .B1(new_n824), .B2(new_n758), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G128), .B2(new_n751), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n764), .C2(new_n1119), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT59), .Z(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n777), .B2(G159), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G33), .B1(new_n779), .B2(G124), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n272), .B1(new_n395), .B2(new_n256), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n322), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n564), .B1(new_n211), .B2(new_n755), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n272), .B1(new_n264), .B2(new_n764), .C1(new_n748), .C2(new_n254), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G116), .C2(new_n771), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n751), .A2(KEYINPUT119), .A3(G107), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT119), .B1(new_n751), .B2(G107), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n778), .A2(new_n810), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n776), .A2(new_n348), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1173), .B(new_n1178), .C1(new_n213), .C2(new_n758), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT58), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1168), .A2(new_n1170), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n746), .B1(new_n1181), .B2(new_n740), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1158), .A2(new_n1159), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT121), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n888), .B2(new_n894), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1157), .B1(new_n876), .B2(G330), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n874), .B1(new_n869), .B2(KEYINPUT40), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1189), .A2(new_n702), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1187), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1189), .B2(new_n702), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n864), .A2(new_n868), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n865), .B1(new_n1194), .B2(new_n841), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1157), .B(G330), .C1(new_n1195), .C2(new_n874), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1193), .A2(new_n1196), .A3(new_n1186), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1184), .B1(new_n1198), .B2(new_n726), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1107), .A2(new_n1101), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1193), .A2(new_n1196), .A3(new_n895), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n895), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(KEYINPUT57), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n677), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1106), .A2(new_n726), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n830), .A2(new_n211), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n759), .A2(G116), .B1(new_n747), .B2(G107), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT122), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G294), .B2(new_n771), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n285), .B1(new_n764), .B2(new_n213), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n752), .A2(new_n810), .B1(new_n755), .B2(new_n254), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G77), .C2(new_n777), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(new_n474), .C2(new_n778), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n755), .A2(new_n322), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n748), .A2(new_n345), .B1(new_n401), .B2(new_n764), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1177), .B(new_n1217), .C1(G128), .C2(new_n779), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n396), .B1(new_n752), .B2(new_n819), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n771), .B2(G132), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n758), .C2(new_n1119), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n746), .B1(new_n1222), .B2(new_n740), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1208), .B(new_n1223), .C1(new_n881), .C2(new_n742), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1207), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT123), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT123), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1207), .A2(new_n1227), .A3(new_n1224), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n902), .A2(new_n650), .A3(new_n1100), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1111), .A2(new_n941), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(G381));
  INV_X1    g1033(.A(new_n1197), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1186), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n726), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1183), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n895), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1193), .A2(new_n1196), .A3(new_n895), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1107), .B2(new_n1101), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n681), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1200), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1242), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1237), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G396), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1045), .A2(new_n1251), .A3(new_n1046), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(G387), .A2(G390), .A3(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G381), .A2(G384), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1253), .A3(new_n1254), .ZN(G407));
  OAI211_X1 g1055(.A(G407), .B(G213), .C1(G343), .C2(new_n1249), .ZN(G409));
  AOI22_X1  g1056(.A1(new_n1192), .A2(new_n1197), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1257), .A2(new_n941), .B1(new_n726), .B2(new_n1241), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1258), .A2(new_n1142), .A3(new_n1116), .A4(new_n1183), .ZN(new_n1259));
  INV_X1    g1059(.A(G213), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(G343), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1259), .B(new_n1262), .C1(new_n1248), .C2(new_n1247), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n681), .B1(new_n1231), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n1111), .C1(new_n1264), .C2(new_n1231), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1229), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1229), .A2(new_n1266), .A3(G384), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(G2897), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1229), .A2(new_n1266), .A3(G384), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n1267), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G375), .A2(G378), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1273), .A2(new_n1267), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1262), .A3(new_n1259), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1116), .A2(new_n1142), .A3(new_n1183), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1241), .A2(new_n726), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1245), .B2(new_n942), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1262), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1276), .A2(new_n1280), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1045), .A2(new_n1251), .A3(new_n1046), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1251), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT125), .A3(new_n1252), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n991), .B1(new_n997), .B2(new_n939), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1074), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1295), .A2(new_n1074), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1293), .B2(new_n1252), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1074), .B1(new_n992), .B2(new_n999), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT126), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1297), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1288), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1203), .B(new_n677), .C1(new_n1257), .C2(KEYINPUT57), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1308), .A2(new_n1199), .B1(new_n1142), .B2(new_n1116), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1284), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT63), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1279), .A2(KEYINPUT124), .A3(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1313), .A2(new_n1302), .A3(new_n1276), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1307), .A2(new_n1316), .ZN(G405));
  NOR2_X1   g1117(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1297), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1304), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1318), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1318), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1303), .A2(new_n1305), .A3(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1250), .A2(new_n1309), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(G402));
endmodule


