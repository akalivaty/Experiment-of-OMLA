//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT67), .Z(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT68), .Z(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT69), .Z(G162));
  OAI211_X1 g056(.A(KEYINPUT4), .B(G138), .C1(new_n460), .C2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(G102), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(KEYINPUT70), .A2(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT70), .A2(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n464), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(new_n462), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(G138), .A3(new_n474), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n484), .B1(new_n494), .B2(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(G88), .B1(new_n510), .B2(G50), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI221_X1 g089(.A(KEYINPUT72), .B1(new_n509), .B2(new_n513), .C1(new_n507), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n505), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(new_n508), .A2(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n509), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n519), .A2(new_n524), .ZN(G168));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n507), .A2(new_n526), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(new_n501), .ZN(new_n532));
  AOI21_X1  g107(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n504), .B1(new_n536), .B2(KEYINPUT73), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n537), .B1(KEYINPUT73), .B2(new_n536), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n530), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n534), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n545), .B(new_n541), .C1(new_n534), .C2(new_n542), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n546), .A3(G651), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT77), .B(G43), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n507), .A2(new_n550), .B1(new_n509), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n547), .B2(new_n548), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n509), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n506), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n563), .A2(new_n565), .B1(new_n508), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n502), .A2(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n504), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(KEYINPUT78), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n571), .B(new_n504), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n566), .B1(new_n570), .B2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(G166), .A2(KEYINPUT79), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n517), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(G303));
  NAND2_X1  g153(.A1(new_n510), .A2(G49), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT80), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n502), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(G87), .A2(new_n508), .B1(new_n581), .B2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n534), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n510), .B2(G48), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n507), .ZN(G305));
  AOI22_X1  g164(.A1(new_n508), .A2(G85), .B1(new_n510), .B2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n504), .B2(new_n591), .ZN(G290));
  XOR2_X1   g167(.A(KEYINPUT83), .B(G66), .Z(new_n593));
  AND2_X1   g168(.A1(new_n593), .A2(new_n502), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT82), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n510), .A2(G54), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n507), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n599), .A2(new_n502), .A3(G92), .A4(new_n506), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n597), .A2(new_n598), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G280));
  AOI21_X1  g186(.A(new_n596), .B1(new_n502), .B2(new_n593), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n598), .B1(new_n612), .B2(new_n504), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n602), .A2(new_n603), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NOR2_X1   g192(.A1(new_n604), .A2(G559), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n556), .B2(G868), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n495), .A2(new_n465), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT13), .Z(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT84), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n463), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n478), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n474), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT85), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n628), .B(new_n635), .C1(new_n626), .C2(new_n625), .ZN(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT86), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT88), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT17), .A3(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n663), .B(new_n664), .C1(new_n662), .C2(new_n658), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n663), .B2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT89), .B(G2100), .Z(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2096), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT90), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n671), .A2(new_n673), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(new_n676), .A3(new_n674), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n681), .C1(new_n676), .C2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT92), .ZN(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n683), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G33), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n463), .A2(G139), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT99), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT25), .Z(new_n697));
  AOI22_X1  g272(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n697), .C1(new_n474), .C2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT100), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n692), .B1(new_n701), .B2(new_n691), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G2072), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT101), .ZN(new_n704));
  INV_X1    g279(.A(G1341), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT96), .B(G16), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G19), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n556), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n704), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n691), .A2(G35), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G162), .B2(new_n691), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT29), .B(G2090), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n691), .A2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n465), .A2(G105), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n463), .A2(G141), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n478), .A2(G129), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT26), .Z(new_n721));
  AND4_X1   g296(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n691), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT27), .B(G1996), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT102), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(new_n691), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n633), .B2(new_n691), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT103), .Z(new_n732));
  NOR2_X1   g307(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n615), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G4), .B2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(G1348), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(G164), .A2(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G27), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G160), .A2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT24), .B2(new_n744), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(G2084), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n733), .A2(new_n738), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n691), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n463), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n478), .A2(G128), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n734), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n734), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1966), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n715), .A2(new_n748), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n706), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n736), .A2(new_n737), .ZN(new_n768));
  AOI21_X1  g343(.A(G2084), .B1(new_n743), .B2(new_n746), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n740), .A2(new_n741), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n734), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n734), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1961), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n710), .A2(new_n705), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G2072), .C2(new_n702), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n711), .A2(new_n762), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n734), .A2(G23), .ZN(new_n778));
  INV_X1    g353(.A(G288), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n734), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT33), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1976), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n707), .A2(G22), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n707), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1971), .Z(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n782), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n463), .A2(G131), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT93), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n478), .A2(G119), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT94), .Z(new_n795));
  INV_X1    g370(.A(G95), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n796), .A2(new_n474), .A3(KEYINPUT95), .ZN(new_n797));
  AOI21_X1  g372(.A(KEYINPUT95), .B1(new_n796), .B2(new_n474), .ZN(new_n798));
  OAI221_X1 g373(.A(G2104), .B1(G107), .B2(new_n474), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G25), .B(new_n800), .S(G29), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT35), .B(G1991), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G24), .B(G290), .S(new_n707), .Z(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT97), .B(G1986), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n790), .A2(new_n791), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n809), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n777), .B1(new_n810), .B2(new_n811), .ZN(G311));
  INV_X1    g387(.A(new_n777), .ZN(new_n813));
  INV_X1    g388(.A(new_n811), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n807), .A2(new_n809), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G150));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT105), .B(G55), .Z(new_n818));
  OAI22_X1  g393(.A1(new_n507), .A2(new_n817), .B1(new_n509), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  INV_X1    g395(.A(G67), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n534), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n504), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n819), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n549), .A2(new_n554), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n549), .B2(new_n554), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n616), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  AOI21_X1  g408(.A(G860), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT106), .Z(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G145));
  NAND2_X1  g415(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n841));
  AND2_X1   g416(.A1(KEYINPUT70), .A2(G114), .ZN(new_n842));
  NOR2_X1   g417(.A1(KEYINPUT70), .A2(G114), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(G126), .B1(new_n460), .B2(new_n461), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n474), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT4), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n496), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n484), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n755), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(new_n722), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n722), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n841), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n800), .B(new_n624), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n841), .A2(new_n855), .A3(new_n852), .A4(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n699), .B(KEYINPUT100), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n463), .A2(G142), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n478), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n474), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n862), .B(new_n867), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n862), .B(new_n867), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n858), .A3(new_n857), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G160), .B(new_n633), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G162), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n871), .ZN(new_n877));
  INV_X1    g452(.A(new_n874), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g454(.A(KEYINPUT108), .B(new_n874), .C1(new_n869), .C2(new_n871), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g457(.A(G288), .B(G305), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n517), .B(G290), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n883), .B(new_n884), .Z(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT42), .Z(new_n886));
  INV_X1    g461(.A(KEYINPUT111), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(G299), .B2(new_n615), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT110), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n569), .B(KEYINPUT78), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n891), .A2(KEYINPUT109), .A3(new_n604), .A4(new_n566), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G299), .A2(new_n615), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n889), .B2(new_n892), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n887), .B1(new_n897), .B2(KEYINPUT41), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  OAI211_X1 g474(.A(KEYINPUT111), .B(new_n899), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n889), .A2(new_n894), .A3(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT41), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n829), .B(new_n619), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n904), .B2(new_n901), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n886), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n886), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G868), .B2(new_n826), .ZN(G295));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n826), .ZN(G331));
  NAND2_X1  g486(.A1(G301), .A2(G168), .ZN(new_n912));
  NAND3_X1  g487(.A1(G286), .A2(new_n530), .A3(new_n538), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n829), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n828), .B2(new_n827), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n898), .A2(new_n900), .A3(new_n918), .A4(new_n902), .ZN(new_n919));
  INV_X1    g494(.A(new_n885), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n901), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n919), .B2(new_n922), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(KEYINPUT43), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n921), .A2(new_n897), .A3(new_n899), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n885), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n901), .B1(new_n921), .B2(new_n899), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n919), .A2(new_n922), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n885), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n928), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n927), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n925), .B2(new_n926), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n934), .A3(new_n928), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n941), .B2(new_n936), .ZN(new_n942));
  AOI211_X1 g517(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n939), .C2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(G397));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n850), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n755), .B(G2067), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n950), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n722), .B(G1996), .ZN(new_n954));
  OAI22_X1  g529(.A1(new_n952), .A2(KEYINPUT113), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(KEYINPUT113), .B2(new_n952), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n800), .B(new_n802), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(G1986), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n950), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n575), .A2(G8), .A3(new_n577), .ZN(new_n961));
  NAND2_X1  g536(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n946), .A2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(new_n949), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n850), .A2(new_n969), .A3(new_n945), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(G2090), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n947), .A2(G1384), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n949), .B1(new_n850), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n948), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT114), .B(G1971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n966), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n965), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(G305), .A2(G1981), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT116), .B(G86), .Z(new_n981));
  NAND2_X1  g556(.A1(new_n508), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n587), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT49), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n946), .A2(new_n949), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n966), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n980), .B(KEYINPUT49), .C1(new_n983), .C2(new_n984), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n989), .B(new_n993), .C1(new_n992), .C2(G288), .ZN(new_n994));
  INV_X1    g569(.A(new_n989), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT52), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n991), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n979), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n970), .A2(KEYINPUT117), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n850), .A2(new_n1001), .A3(new_n969), .A4(new_n945), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1000), .A2(new_n967), .A3(new_n968), .A4(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1003), .A2(G2090), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n966), .B1(new_n1004), .B2(new_n977), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n965), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2084), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n967), .A2(new_n1009), .A3(new_n968), .A4(new_n970), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1966), .B1(new_n948), .B2(new_n974), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(KEYINPUT118), .ZN(new_n1012));
  INV_X1    g587(.A(G1966), .ZN(new_n1013));
  INV_X1    g588(.A(new_n973), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n968), .B1(G164), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n850), .B2(new_n945), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT118), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(G8), .B(G286), .C1(new_n1012), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1027), .A2(G168), .A3(new_n1017), .A4(new_n1010), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(KEYINPUT124), .B2(KEYINPUT51), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1024), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1020), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1030), .A3(new_n1024), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT125), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1023), .ZN(new_n1036));
  AND4_X1   g611(.A1(KEYINPUT125), .A2(new_n1036), .A3(new_n1033), .A4(new_n1019), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT62), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1033), .A3(new_n1019), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1032), .A2(KEYINPUT125), .A3(new_n1033), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n975), .B2(G2078), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT53), .A3(new_n741), .ZN(new_n1048));
  INV_X1    g623(.A(G1961), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n971), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT126), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1038), .A2(new_n1044), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1051), .A2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1052), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1056), .A2(KEYINPUT127), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OR3_X1    g635(.A1(new_n1051), .A2(G171), .A3(new_n1059), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1054), .A2(new_n1056), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n988), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G2067), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n971), .A2(new_n737), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n604), .B(KEYINPUT123), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(KEYINPUT60), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1066), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(new_n1064), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1070), .A2(new_n1069), .A3(new_n1064), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n615), .A2(KEYINPUT123), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1068), .B(new_n1071), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT61), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1003), .A2(new_n766), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G299), .A2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT57), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1047), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1079), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1075), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1996), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1047), .A2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n1063), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n555), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1076), .A2(new_n1081), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1079), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1082), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1074), .A2(new_n1085), .A3(new_n1092), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n604), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1082), .B1(new_n1098), .B2(new_n1084), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1062), .B(new_n1100), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1008), .B1(new_n1055), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n991), .A2(new_n992), .A3(new_n779), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n995), .B1(new_n1103), .B2(new_n980), .ZN(new_n1104));
  INV_X1    g679(.A(new_n979), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n998), .ZN(new_n1106));
  OAI211_X1 g681(.A(G8), .B(G168), .C1(new_n1012), .C2(new_n1018), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT119), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT63), .A3(new_n979), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n998), .B1(new_n965), .B2(new_n978), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1007), .B2(new_n1108), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1106), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n960), .B1(new_n1102), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n950), .A2(new_n1086), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT46), .ZN(new_n1119));
  INV_X1    g694(.A(new_n722), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n951), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1118), .A2(new_n1119), .B1(new_n950), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1119), .B2(new_n1118), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT47), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n953), .A2(G1986), .A3(G290), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT48), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n958), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n802), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n800), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n956), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n755), .A2(G2067), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n953), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1117), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(G319), .ZN(new_n1136));
  NOR4_X1   g710(.A1(G401), .A2(new_n1136), .A3(G227), .A4(G229), .ZN(new_n1137));
  NAND3_X1  g711(.A1(new_n881), .A2(new_n941), .A3(new_n1137), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


