

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731;

  XNOR2_X1 U366 ( .A(n553), .B(n552), .ZN(n585) );
  OR2_X1 U367 ( .A1(n374), .A2(n471), .ZN(n474) );
  INV_X2 U368 ( .A(G953), .ZN(n718) );
  NOR2_X1 U369 ( .A1(n527), .A2(n505), .ZN(n636) );
  XNOR2_X2 U370 ( .A(n591), .B(n590), .ZN(n699) );
  NAND2_X1 U371 ( .A1(n650), .A2(n649), .ZN(n574) );
  NOR2_X1 U372 ( .A1(n574), .A2(n582), .ZN(n559) );
  AND2_X1 U373 ( .A1(n614), .A2(n613), .ZN(n616) );
  AND2_X1 U374 ( .A1(n619), .A2(n613), .ZN(n621) );
  NOR2_X1 U375 ( .A1(n527), .A2(n680), .ZN(n529) );
  XNOR2_X1 U376 ( .A(n526), .B(n525), .ZN(n680) );
  AND2_X1 U377 ( .A1(n666), .A2(n375), .ZN(n526) );
  OR2_X1 U378 ( .A1(n523), .A2(n496), .ZN(n519) );
  NOR2_X1 U379 ( .A1(n669), .A2(n502), .ZN(n375) );
  XNOR2_X1 U380 ( .A(n422), .B(n421), .ZN(n523) );
  XNOR2_X1 U381 ( .A(n419), .B(n418), .ZN(n595) );
  XNOR2_X1 U382 ( .A(n379), .B(n378), .ZN(n419) );
  XNOR2_X1 U383 ( .A(n417), .B(n349), .ZN(n379) );
  XNOR2_X1 U384 ( .A(n465), .B(G134), .ZN(n444) );
  XNOR2_X1 U385 ( .A(KEYINPUT72), .B(G131), .ZN(n443) );
  NOR2_X4 U386 ( .A1(n647), .A2(n594), .ZN(n688) );
  XNOR2_X2 U387 ( .A(n593), .B(n592), .ZN(n647) );
  XNOR2_X1 U388 ( .A(n354), .B(n353), .ZN(n394) );
  XNOR2_X1 U389 ( .A(n713), .B(n445), .ZN(n485) );
  INV_X1 U390 ( .A(G146), .ZN(n445) );
  XNOR2_X1 U391 ( .A(n411), .B(n410), .ZN(n522) );
  XNOR2_X1 U392 ( .A(n409), .B(n408), .ZN(n410) );
  BUF_X1 U393 ( .A(n498), .Z(n573) );
  XNOR2_X1 U394 ( .A(n370), .B(n369), .ZN(n368) );
  INV_X1 U395 ( .A(KEYINPUT28), .ZN(n369) );
  NAND2_X1 U396 ( .A1(n499), .A2(n371), .ZN(n370) );
  NOR2_X1 U397 ( .A1(KEYINPUT47), .A2(n579), .ZN(n497) );
  XNOR2_X1 U398 ( .A(n452), .B(n451), .ZN(n498) );
  NAND2_X1 U399 ( .A1(n645), .A2(n390), .ZN(n387) );
  INV_X1 U400 ( .A(KEYINPUT87), .ZN(n390) );
  INV_X1 U401 ( .A(n643), .ZN(n392) );
  NAND2_X1 U402 ( .A1(n394), .A2(n347), .ZN(n388) );
  XNOR2_X1 U403 ( .A(n444), .B(n373), .ZN(n713) );
  INV_X1 U404 ( .A(n443), .ZN(n373) );
  NOR2_X1 U405 ( .A1(n726), .A2(n571), .ZN(n572) );
  XNOR2_X1 U406 ( .A(n377), .B(KEYINPUT71), .ZN(n412) );
  INV_X1 U407 ( .A(KEYINPUT10), .ZN(n377) );
  XNOR2_X1 U408 ( .A(G137), .B(G140), .ZN(n424) );
  XNOR2_X1 U409 ( .A(n364), .B(G101), .ZN(n478) );
  INV_X1 U410 ( .A(KEYINPUT4), .ZN(n364) );
  INV_X1 U411 ( .A(G107), .ZN(n476) );
  XNOR2_X1 U412 ( .A(n363), .B(n491), .ZN(n516) );
  NOR2_X1 U413 ( .A1(n362), .A2(n361), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n420), .B(G475), .ZN(n421) );
  NOR2_X1 U415 ( .A1(G902), .A2(n595), .ZN(n422) );
  XNOR2_X1 U416 ( .A(n433), .B(n432), .ZN(n500) );
  XNOR2_X1 U417 ( .A(n456), .B(G104), .ZN(n480) );
  XNOR2_X1 U418 ( .A(KEYINPUT91), .B(G110), .ZN(n456) );
  XNOR2_X1 U419 ( .A(KEYINPUT3), .B(G119), .ZN(n704) );
  XNOR2_X1 U420 ( .A(n382), .B(n381), .ZN(n380) );
  XNOR2_X1 U421 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U422 ( .A(KEYINPUT94), .B(KEYINPUT85), .ZN(n382) );
  NAND2_X1 U423 ( .A1(n455), .A2(n372), .ZN(n535) );
  XNOR2_X1 U424 ( .A(n504), .B(n503), .ZN(n548) );
  OR2_X1 U425 ( .A1(n538), .A2(n502), .ZN(n504) );
  INV_X1 U426 ( .A(G469), .ZN(n400) );
  NOR2_X1 U427 ( .A1(G902), .A2(n604), .ZN(n486) );
  XNOR2_X1 U428 ( .A(n407), .B(n406), .ZN(n690) );
  XNOR2_X1 U429 ( .A(n670), .B(KEYINPUT84), .ZN(n579) );
  AND2_X1 U430 ( .A1(n519), .A2(n542), .ZN(n670) );
  NOR2_X1 U431 ( .A1(n489), .A2(n490), .ZN(n362) );
  NOR2_X1 U432 ( .A1(n667), .A2(n490), .ZN(n361) );
  NAND2_X1 U433 ( .A1(n358), .A2(n356), .ZN(n355) );
  AND2_X1 U434 ( .A1(n654), .A2(n346), .ZN(n399) );
  XNOR2_X1 U435 ( .A(G128), .B(G110), .ZN(n384) );
  XNOR2_X1 U436 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n385) );
  XNOR2_X1 U437 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n381) );
  XNOR2_X1 U438 ( .A(G143), .B(G140), .ZN(n416) );
  XNOR2_X1 U439 ( .A(n415), .B(n425), .ZN(n378) );
  XOR2_X1 U440 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n414) );
  XNOR2_X1 U441 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n427) );
  AND2_X1 U442 ( .A1(n500), .A2(n346), .ZN(n371) );
  NOR2_X1 U443 ( .A1(n543), .A2(n498), .ZN(n499) );
  XNOR2_X1 U444 ( .A(n485), .B(n365), .ZN(n611) );
  XNOR2_X1 U445 ( .A(n366), .B(n468), .ZN(n365) );
  XNOR2_X1 U446 ( .A(n448), .B(n348), .ZN(n366) );
  NOR2_X1 U447 ( .A1(n394), .A2(KEYINPUT87), .ZN(n391) );
  NAND2_X1 U448 ( .A1(n388), .A2(n386), .ZN(n389) );
  AND2_X1 U449 ( .A1(n387), .A2(n392), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n484), .B(n485), .ZN(n604) );
  NOR2_X1 U451 ( .A1(n673), .A2(n560), .ZN(n561) );
  NAND2_X1 U452 ( .A1(n523), .A2(n496), .ZN(n542) );
  INV_X1 U453 ( .A(G101), .ZN(n705) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n696) );
  XNOR2_X1 U455 ( .A(n426), .B(G119), .ZN(n395) );
  NOR2_X1 U456 ( .A1(n535), .A2(n538), .ZN(n475) );
  INV_X1 U457 ( .A(KEYINPUT104), .ZN(n492) );
  INV_X1 U458 ( .A(n542), .ZN(n639) );
  NAND2_X1 U459 ( .A1(n345), .A2(n356), .ZN(n576) );
  XNOR2_X1 U460 ( .A(n690), .B(n689), .ZN(n691) );
  INV_X1 U461 ( .A(n645), .ZN(n393) );
  NOR2_X2 U462 ( .A1(n391), .A2(n389), .ZN(n716) );
  XOR2_X1 U463 ( .A(n383), .B(n380), .Z(n344) );
  AND2_X1 U464 ( .A1(n501), .A2(n654), .ZN(n345) );
  AND2_X1 U465 ( .A1(n440), .A2(n648), .ZN(n346) );
  AND2_X1 U466 ( .A1(n393), .A2(KEYINPUT87), .ZN(n347) );
  AND2_X1 U467 ( .A1(n449), .A2(G210), .ZN(n348) );
  AND2_X1 U468 ( .A1(G214), .A2(n449), .ZN(n349) );
  OR2_X1 U469 ( .A1(n543), .A2(n454), .ZN(n350) );
  XOR2_X1 U470 ( .A(n374), .B(n617), .Z(n351) );
  XNOR2_X1 U471 ( .A(KEYINPUT62), .B(n611), .ZN(n352) );
  XOR2_X1 U472 ( .A(KEYINPUT48), .B(KEYINPUT74), .Z(n353) );
  NAND2_X1 U473 ( .A1(n533), .A2(n534), .ZN(n354) );
  NOR2_X1 U474 ( .A1(n355), .A2(n398), .ZN(n357) );
  INV_X1 U475 ( .A(n500), .ZN(n356) );
  NAND2_X1 U476 ( .A1(n360), .A2(n357), .ZN(n363) );
  NAND2_X1 U477 ( .A1(n489), .A2(n359), .ZN(n358) );
  AND2_X1 U478 ( .A1(n667), .A2(n490), .ZN(n359) );
  NAND2_X1 U479 ( .A1(n727), .A2(n367), .ZN(n532) );
  XNOR2_X1 U480 ( .A(n367), .B(G137), .ZN(G39) );
  XNOR2_X1 U481 ( .A(n530), .B(KEYINPUT106), .ZN(n367) );
  NAND2_X1 U482 ( .A1(n368), .A2(n501), .ZN(n527) );
  NOR2_X1 U483 ( .A1(n582), .A2(n350), .ZN(n372) );
  XNOR2_X2 U484 ( .A(G143), .B(G128), .ZN(n465) );
  XNOR2_X1 U485 ( .A(n707), .B(n470), .ZN(n374) );
  NAND2_X1 U486 ( .A1(n666), .A2(n667), .ZN(n376) );
  NOR2_X1 U487 ( .A1(n670), .A2(n376), .ZN(n671) );
  NOR2_X1 U488 ( .A1(n729), .A2(n513), .ZN(n534) );
  NOR2_X1 U489 ( .A1(n696), .A2(G902), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n712), .B(n344), .ZN(n396) );
  XNOR2_X1 U491 ( .A(n425), .B(n397), .ZN(n712) );
  INV_X1 U492 ( .A(n481), .ZN(n397) );
  NAND2_X1 U493 ( .A1(n501), .A2(n399), .ZN(n398) );
  XNOR2_X2 U494 ( .A(n486), .B(n400), .ZN(n501) );
  NOR2_X1 U495 ( .A1(n500), .A2(n543), .ZN(n650) );
  NOR2_X1 U496 ( .A1(n541), .A2(n519), .ZN(n521) );
  XNOR2_X2 U497 ( .A(n501), .B(KEYINPUT1), .ZN(n649) );
  XNOR2_X1 U498 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U499 ( .A(n479), .B(n478), .ZN(n483) );
  INV_X1 U500 ( .A(KEYINPUT30), .ZN(n490) );
  INV_X1 U501 ( .A(KEYINPUT100), .ZN(n408) );
  XNOR2_X1 U502 ( .A(n443), .B(KEYINPUT98), .ZN(n418) );
  NOR2_X1 U503 ( .A1(n516), .A2(n524), .ZN(n518) );
  INV_X1 U504 ( .A(KEYINPUT81), .ZN(n491) );
  XNOR2_X1 U505 ( .A(n444), .B(n405), .ZN(n406) );
  INV_X1 U506 ( .A(KEYINPUT66), .ZN(n555) );
  XNOR2_X1 U507 ( .A(n556), .B(n555), .ZN(n557) );
  INV_X1 U508 ( .A(n698), .ZN(n613) );
  XNOR2_X1 U509 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U510 ( .A1(G234), .A2(n718), .ZN(n402) );
  XOR2_X1 U511 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n401) );
  XNOR2_X1 U512 ( .A(n402), .B(n401), .ZN(n423) );
  NAND2_X1 U513 ( .A1(G217), .A2(n423), .ZN(n404) );
  XNOR2_X1 U514 ( .A(G116), .B(G107), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT7), .ZN(n403) );
  XNOR2_X1 U516 ( .A(n404), .B(n403), .ZN(n407) );
  XNOR2_X1 U517 ( .A(G122), .B(KEYINPUT9), .ZN(n405) );
  NOR2_X1 U518 ( .A1(G902), .A2(n690), .ZN(n411) );
  INV_X1 U519 ( .A(G478), .ZN(n409) );
  INV_X1 U520 ( .A(n522), .ZN(n496) );
  XNOR2_X2 U521 ( .A(G146), .B(G125), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n412), .B(n464), .ZN(n425) );
  XNOR2_X1 U523 ( .A(G104), .B(KEYINPUT11), .ZN(n413) );
  XNOR2_X1 U524 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U525 ( .A1(G953), .A2(G237), .ZN(n449) );
  XNOR2_X1 U526 ( .A(G122), .B(G113), .ZN(n457) );
  XNOR2_X1 U527 ( .A(n457), .B(n416), .ZN(n417) );
  XNOR2_X1 U528 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n420) );
  XOR2_X1 U529 ( .A(KEYINPUT102), .B(n519), .Z(n623) );
  NAND2_X1 U530 ( .A1(G221), .A2(n423), .ZN(n426) );
  XNOR2_X1 U531 ( .A(n424), .B(KEYINPUT73), .ZN(n481) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(KEYINPUT82), .Z(n430) );
  XNOR2_X1 U533 ( .A(n427), .B(G902), .ZN(n594) );
  NAND2_X1 U534 ( .A1(n594), .A2(G234), .ZN(n428) );
  XNOR2_X1 U535 ( .A(KEYINPUT20), .B(n428), .ZN(n441) );
  NAND2_X1 U536 ( .A1(n441), .A2(G217), .ZN(n429) );
  XNOR2_X1 U537 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U538 ( .A(n431), .B(KEYINPUT96), .ZN(n432) );
  INV_X1 U539 ( .A(n356), .ZN(n581) );
  AND2_X1 U540 ( .A1(n623), .A2(n581), .ZN(n455) );
  INV_X1 U541 ( .A(G902), .ZN(n450) );
  INV_X1 U542 ( .A(G237), .ZN(n434) );
  NAND2_X1 U543 ( .A1(n450), .A2(n434), .ZN(n472) );
  NAND2_X1 U544 ( .A1(n472), .A2(G214), .ZN(n667) );
  NOR2_X1 U545 ( .A1(G900), .A2(n718), .ZN(n435) );
  NAND2_X1 U546 ( .A1(n435), .A2(G902), .ZN(n436) );
  NAND2_X1 U547 ( .A1(G952), .A2(n718), .ZN(n544) );
  NAND2_X1 U548 ( .A1(n436), .A2(n544), .ZN(n440) );
  XOR2_X1 U549 ( .A(KEYINPUT92), .B(KEYINPUT14), .Z(n438) );
  NAND2_X1 U550 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U551 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U552 ( .A(n439), .B(KEYINPUT79), .ZN(n648) );
  NAND2_X1 U553 ( .A1(n667), .A2(n346), .ZN(n454) );
  AND2_X1 U554 ( .A1(n441), .A2(G221), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n442), .B(KEYINPUT21), .ZN(n654) );
  INV_X1 U556 ( .A(n654), .ZN(n543) );
  XNOR2_X1 U557 ( .A(n478), .B(n704), .ZN(n468) );
  XOR2_X1 U558 ( .A(KEYINPUT5), .B(G113), .Z(n447) );
  XNOR2_X1 U559 ( .A(G137), .B(G116), .ZN(n446) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n448) );
  NAND2_X1 U561 ( .A1(n611), .A2(n450), .ZN(n452) );
  INV_X1 U562 ( .A(G472), .ZN(n451) );
  INV_X1 U563 ( .A(KEYINPUT6), .ZN(n453) );
  XNOR2_X1 U564 ( .A(n573), .B(n453), .ZN(n582) );
  XNOR2_X1 U565 ( .A(n480), .B(n457), .ZN(n461) );
  XNOR2_X1 U566 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n461), .B(n460), .ZN(n707) );
  XNOR2_X1 U569 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n463) );
  NAND2_X1 U570 ( .A1(n718), .A2(G224), .ZN(n462) );
  XNOR2_X1 U571 ( .A(n463), .B(n462), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U573 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U575 ( .A(n594), .ZN(n471) );
  NAND2_X1 U576 ( .A1(n472), .A2(G210), .ZN(n473) );
  XNOR2_X2 U577 ( .A(n474), .B(n473), .ZN(n538) );
  XNOR2_X1 U578 ( .A(n475), .B(KEYINPUT36), .ZN(n487) );
  NAND2_X1 U579 ( .A1(G227), .A2(n718), .ZN(n477) );
  XNOR2_X1 U580 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U581 ( .A(n483), .B(n482), .Z(n484) );
  XOR2_X1 U582 ( .A(KEYINPUT89), .B(n649), .Z(n566) );
  NAND2_X1 U583 ( .A1(n487), .A2(n566), .ZN(n488) );
  XNOR2_X1 U584 ( .A(n488), .B(KEYINPUT107), .ZN(n729) );
  NOR2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n562) );
  INV_X1 U586 ( .A(n562), .ZN(n495) );
  INV_X1 U587 ( .A(n498), .ZN(n489) );
  NOR2_X1 U588 ( .A1(n516), .A2(n538), .ZN(n493) );
  XNOR2_X1 U589 ( .A(n493), .B(n492), .ZN(n494) );
  NOR2_X1 U590 ( .A1(n495), .A2(n494), .ZN(n635) );
  XNOR2_X1 U591 ( .A(KEYINPUT78), .B(n497), .ZN(n506) );
  INV_X1 U592 ( .A(n667), .ZN(n502) );
  XNOR2_X1 U593 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n503) );
  INV_X1 U594 ( .A(n548), .ZN(n505) );
  NAND2_X1 U595 ( .A1(n506), .A2(n636), .ZN(n510) );
  INV_X1 U596 ( .A(n670), .ZN(n507) );
  NAND2_X1 U597 ( .A1(n636), .A2(n507), .ZN(n508) );
  NAND2_X1 U598 ( .A1(n508), .A2(KEYINPUT47), .ZN(n509) );
  NAND2_X1 U599 ( .A1(n510), .A2(n509), .ZN(n511) );
  NOR2_X1 U600 ( .A1(n635), .A2(n511), .ZN(n512) );
  XNOR2_X1 U601 ( .A(n512), .B(KEYINPUT77), .ZN(n513) );
  INV_X1 U602 ( .A(KEYINPUT80), .ZN(n514) );
  XNOR2_X1 U603 ( .A(n514), .B(KEYINPUT38), .ZN(n515) );
  XNOR2_X1 U604 ( .A(n538), .B(n515), .ZN(n524) );
  XNOR2_X1 U605 ( .A(KEYINPUT39), .B(KEYINPUT88), .ZN(n517) );
  XNOR2_X1 U606 ( .A(n518), .B(n517), .ZN(n541) );
  INV_X1 U607 ( .A(KEYINPUT40), .ZN(n520) );
  XNOR2_X1 U608 ( .A(n521), .B(n520), .ZN(n727) );
  NAND2_X1 U609 ( .A1(n523), .A2(n522), .ZN(n669) );
  INV_X1 U610 ( .A(n524), .ZN(n666) );
  XOR2_X1 U611 ( .A(KEYINPUT41), .B(KEYINPUT105), .Z(n525) );
  INV_X1 U612 ( .A(KEYINPUT42), .ZN(n528) );
  XNOR2_X1 U613 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U614 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n531) );
  XNOR2_X1 U615 ( .A(n532), .B(n531), .ZN(n533) );
  NOR2_X1 U616 ( .A1(n535), .A2(n649), .ZN(n536) );
  XNOR2_X1 U617 ( .A(n536), .B(KEYINPUT103), .ZN(n537) );
  XOR2_X1 U618 ( .A(KEYINPUT43), .B(n537), .Z(n540) );
  INV_X1 U619 ( .A(n538), .ZN(n539) );
  NOR2_X1 U620 ( .A1(n540), .A2(n539), .ZN(n645) );
  NOR2_X1 U621 ( .A1(n541), .A2(n542), .ZN(n643) );
  NOR2_X1 U622 ( .A1(n669), .A2(n543), .ZN(n551) );
  NOR2_X1 U623 ( .A1(G898), .A2(n718), .ZN(n709) );
  NAND2_X1 U624 ( .A1(G902), .A2(n709), .ZN(n545) );
  NAND2_X1 U625 ( .A1(n545), .A2(n544), .ZN(n546) );
  AND2_X1 U626 ( .A1(n648), .A2(n546), .ZN(n547) );
  NAND2_X1 U627 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U628 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n549) );
  XNOR2_X2 U629 ( .A(n550), .B(n549), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n551), .A2(n577), .ZN(n553) );
  XNOR2_X1 U631 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n552) );
  INV_X1 U632 ( .A(n573), .ZN(n657) );
  NOR2_X1 U633 ( .A1(n649), .A2(n657), .ZN(n554) );
  NAND2_X1 U634 ( .A1(n585), .A2(n554), .ZN(n556) );
  NAND2_X1 U635 ( .A1(n557), .A2(n581), .ZN(n558) );
  XNOR2_X1 U636 ( .A(n558), .B(KEYINPUT101), .ZN(n726) );
  XNOR2_X1 U637 ( .A(n559), .B(KEYINPUT33), .ZN(n673) );
  INV_X1 U638 ( .A(n577), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n561), .B(KEYINPUT34), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U641 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n564) );
  XNOR2_X1 U642 ( .A(n565), .B(n564), .ZN(n725) );
  INV_X1 U643 ( .A(n566), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n567) );
  NOR2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U646 ( .A1(n569), .A2(n585), .ZN(n570) );
  XNOR2_X1 U647 ( .A(n570), .B(KEYINPUT32), .ZN(n610) );
  NAND2_X1 U648 ( .A1(n725), .A2(n610), .ZN(n571) );
  XNOR2_X1 U649 ( .A(n572), .B(KEYINPUT44), .ZN(n588) );
  NOR2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n663) );
  NAND2_X1 U651 ( .A1(n663), .A2(n577), .ZN(n575) );
  XNOR2_X1 U652 ( .A(n575), .B(KEYINPUT31), .ZN(n640) );
  NOR2_X1 U653 ( .A1(n576), .A2(n657), .ZN(n578) );
  AND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n626) );
  NOR2_X1 U655 ( .A1(n640), .A2(n626), .ZN(n580) );
  NOR2_X1 U656 ( .A1(n580), .A2(n579), .ZN(n586) );
  NOR2_X1 U657 ( .A1(n649), .A2(n581), .ZN(n583) );
  AND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n622) );
  NOR2_X1 U660 ( .A1(n586), .A2(n622), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT86), .B(KEYINPUT45), .Z(n589) );
  XNOR2_X1 U663 ( .A(n589), .B(KEYINPUT65), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n716), .A2(n699), .ZN(n593) );
  INV_X1 U665 ( .A(KEYINPUT2), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n688), .A2(G475), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT67), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n599), .B(n598), .ZN(n601) );
  INV_X1 U671 ( .A(G952), .ZN(n600) );
  AND2_X1 U672 ( .A1(n600), .A2(G953), .ZN(n698) );
  NOR2_X2 U673 ( .A1(n601), .A2(n698), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U675 ( .A1(n688), .A2(G469), .ZN(n606) );
  XOR2_X1 U676 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n603) );
  XNOR2_X1 U677 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n607) );
  INV_X1 U679 ( .A(n607), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n608), .A2(n613), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT123), .ZN(G54) );
  XNOR2_X1 U682 ( .A(n610), .B(G119), .ZN(G21) );
  NAND2_X1 U683 ( .A1(n688), .A2(G472), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(n352), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT108), .B(KEYINPUT63), .Z(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(G57) );
  NAND2_X1 U687 ( .A1(n688), .A2(G210), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n351), .ZN(n619) );
  XNOR2_X1 U690 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G51) );
  XOR2_X1 U692 ( .A(G101), .B(n622), .Z(G3) );
  XOR2_X1 U693 ( .A(G104), .B(KEYINPUT109), .Z(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n623), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  NAND2_X1 U697 ( .A1(n626), .A2(n639), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U699 ( .A(G107), .B(n629), .ZN(G9) );
  XOR2_X1 U700 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n631) );
  XNOR2_X1 U701 ( .A(G128), .B(KEYINPUT111), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U703 ( .A(KEYINPUT110), .B(n632), .Z(n634) );
  NAND2_X1 U704 ( .A1(n636), .A2(n639), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G30) );
  XOR2_X1 U706 ( .A(G143), .B(n635), .Z(G45) );
  NAND2_X1 U707 ( .A1(n623), .A2(n636), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(G146), .ZN(G48) );
  NAND2_X1 U709 ( .A1(n623), .A2(n640), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(G113), .ZN(G15) );
  XOR2_X1 U711 ( .A(G116), .B(KEYINPUT113), .Z(n642) );
  NAND2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G18) );
  XNOR2_X1 U714 ( .A(G134), .B(n643), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n644), .B(KEYINPUT115), .ZN(G36) );
  XOR2_X1 U716 ( .A(G140), .B(n645), .Z(n646) );
  XNOR2_X1 U717 ( .A(KEYINPUT116), .B(n646), .ZN(G42) );
  INV_X1 U718 ( .A(n647), .ZN(n685) );
  NAND2_X1 U719 ( .A1(G952), .A2(n648), .ZN(n679) );
  NOR2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U721 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U723 ( .A(KEYINPUT118), .B(n653), .Z(n660) );
  NOR2_X1 U724 ( .A1(n356), .A2(n654), .ZN(n655) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(n655), .Z(n656) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(KEYINPUT117), .B(n658), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT120), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U731 ( .A(KEYINPUT51), .B(n664), .Z(n665) );
  NOR2_X1 U732 ( .A1(n680), .A2(n665), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U738 ( .A(n677), .B(KEYINPUT52), .ZN(n678) );
  NOR2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n682) );
  NOR2_X1 U740 ( .A1(n673), .A2(n680), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U742 ( .A1(n683), .A2(n718), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U744 ( .A(KEYINPUT53), .B(n686), .Z(n687) );
  XNOR2_X1 U745 ( .A(KEYINPUT121), .B(n687), .ZN(G75) );
  BUF_X1 U746 ( .A(n688), .Z(n694) );
  NAND2_X1 U747 ( .A1(n694), .A2(G478), .ZN(n692) );
  INV_X1 U748 ( .A(KEYINPUT125), .ZN(n689) );
  NOR2_X1 U749 ( .A1(n698), .A2(n693), .ZN(G63) );
  NAND2_X1 U750 ( .A1(n694), .A2(G217), .ZN(n695) );
  XNOR2_X1 U751 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U752 ( .A1(n698), .A2(n697), .ZN(G66) );
  NAND2_X1 U753 ( .A1(n699), .A2(n718), .ZN(n703) );
  NAND2_X1 U754 ( .A1(G953), .A2(G224), .ZN(n700) );
  XNOR2_X1 U755 ( .A(KEYINPUT61), .B(n700), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n701), .A2(G898), .ZN(n702) );
  NAND2_X1 U757 ( .A1(n703), .A2(n702), .ZN(n711) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(G69) );
  XNOR2_X1 U762 ( .A(n712), .B(KEYINPUT126), .ZN(n715) );
  XNOR2_X1 U763 ( .A(n713), .B(KEYINPUT4), .ZN(n714) );
  XOR2_X1 U764 ( .A(n715), .B(n714), .Z(n720) );
  INV_X1 U765 ( .A(n720), .ZN(n717) );
  XOR2_X1 U766 ( .A(n717), .B(n716), .Z(n719) );
  NAND2_X1 U767 ( .A1(n719), .A2(n718), .ZN(n724) );
  XOR2_X1 U768 ( .A(G227), .B(n720), .Z(n721) );
  NAND2_X1 U769 ( .A1(n721), .A2(G900), .ZN(n722) );
  NAND2_X1 U770 ( .A1(n722), .A2(G953), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n724), .A2(n723), .ZN(G72) );
  XNOR2_X1 U772 ( .A(G122), .B(n725), .ZN(G24) );
  XOR2_X1 U773 ( .A(G110), .B(n726), .Z(G12) );
  XOR2_X1 U774 ( .A(n727), .B(G131), .Z(n728) );
  XNOR2_X1 U775 ( .A(KEYINPUT127), .B(n728), .ZN(G33) );
  XNOR2_X1 U776 ( .A(n729), .B(KEYINPUT114), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT37), .ZN(n731) );
  XNOR2_X1 U778 ( .A(G125), .B(n731), .ZN(G27) );
endmodule

