//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G22gat), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT31), .ZN(new_n206));
  INV_X1    g005(.A(G228gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT79), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G162gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n213), .A3(G155gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G155gat), .B(G162gat), .Z(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n222));
  OAI21_X1  g021(.A(G141gat), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n218), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n214), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n217), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(KEYINPUT77), .ZN(new_n227));
  XNOR2_X1  g026(.A(G155gat), .B(G162gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G141gat), .B(G148gat), .Z(new_n232));
  INV_X1    g031(.A(G155gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT2), .B1(new_n233), .B2(new_n210), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n226), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n238), .B2(new_n240), .ZN(new_n243));
  XNOR2_X1  g042(.A(G197gat), .B(G204gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n245));
  INV_X1    g044(.A(G211gat), .ZN(new_n246));
  INV_X1    g045(.A(G218gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G211gat), .B(G218gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT75), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n242), .A2(new_n243), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n240), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n237), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n226), .A2(new_n236), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n209), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n251), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n240), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n209), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n257), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n206), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(KEYINPUT83), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n261), .A3(new_n241), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n268), .B2(new_n257), .ZN(new_n269));
  INV_X1    g068(.A(new_n265), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n269), .A2(KEYINPUT31), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n205), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n259), .A2(new_n206), .A3(new_n265), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT31), .B1(new_n269), .B2(new_n270), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n204), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277));
  INV_X1    g076(.A(G113gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(G120gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(G113gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(G113gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(G120gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT68), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT69), .B(G113gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(new_n280), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n288), .A2(new_n283), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n287), .A2(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  AND2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(KEYINPUT24), .ZN(new_n296));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT64), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n301), .A3(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n296), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT25), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n310), .A2(KEYINPUT65), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(KEYINPUT65), .ZN(new_n312));
  OAI211_X1 g111(.A(KEYINPUT23), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n303), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT26), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n306), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n324), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n319), .A2(new_n297), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n305), .A2(new_n307), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n297), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g133(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n296), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n328), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n293), .B1(new_n327), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n286), .A2(new_n283), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT68), .B1(new_n284), .B2(new_n285), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n289), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n292), .A2(new_n291), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  XOR2_X1   g147(.A(KEYINPUT67), .B(KEYINPUT24), .Z(new_n349));
  AND3_X1   g148(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT25), .B1(new_n353), .B2(new_n331), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n346), .A2(new_n354), .A3(new_n314), .A4(new_n326), .ZN(new_n355));
  INV_X1    g154(.A(G227gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(new_n208), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT71), .ZN(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G71gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(G99gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n358), .A2(new_n367), .A3(KEYINPUT32), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n360), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n363), .A2(new_n365), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n341), .A2(new_n355), .ZN(new_n373));
  INV_X1    g172(.A(new_n357), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n372), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n369), .A2(new_n372), .A3(KEYINPUT73), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n372), .ZN(new_n385));
  INV_X1    g184(.A(new_n380), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n276), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n354), .A2(new_n314), .A3(new_n326), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(new_n240), .B1(G226gat), .B2(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n327), .A2(new_n340), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n252), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n392), .B2(KEYINPUT29), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(G226gat), .A3(G233gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n261), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  INV_X1    g199(.A(G64gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G92gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n389), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI211_X1 g206(.A(KEYINPUT30), .B(new_n404), .C1(new_n395), .C2(new_n398), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n405), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT76), .B1(new_n399), .B2(new_n405), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n407), .A2(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G57gat), .ZN(new_n415));
  INV_X1    g214(.A(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n293), .A2(new_n226), .A3(new_n236), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT82), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n293), .A2(new_n226), .A3(new_n420), .A4(new_n236), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(KEYINPUT4), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n423));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT1), .B1(new_n424), .B2(KEYINPUT68), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n288), .B1(new_n425), .B2(new_n282), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n288), .A2(new_n283), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n429));
  OAI21_X1  g228(.A(G120gat), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n284), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT81), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n344), .A2(new_n433), .A3(new_n345), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n423), .A2(new_n435), .A3(new_n238), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT5), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n422), .A2(new_n436), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n293), .A2(new_n226), .A3(KEYINPUT4), .A4(new_n236), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n443), .A2(new_n439), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT4), .B1(new_n419), .B2(new_n421), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n419), .A2(new_n421), .B1(new_n256), .B2(new_n435), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT5), .B1(new_n448), .B2(new_n439), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n417), .B(new_n442), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n214), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT80), .B1(new_n214), .B2(KEYINPUT2), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n455), .A2(new_n224), .B1(new_n235), .B2(new_n231), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n420), .B1(new_n456), .B2(new_n293), .ZN(new_n457));
  INV_X1    g256(.A(new_n421), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n437), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n444), .A3(new_n436), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n435), .A2(new_n256), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n457), .B2(new_n458), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n440), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(KEYINPUT5), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n417), .B1(new_n464), .B2(new_n442), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n452), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n442), .B1(new_n447), .B2(new_n449), .ZN(new_n467));
  INV_X1    g266(.A(new_n417), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n412), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n388), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n383), .A2(new_n384), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT74), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n358), .A2(new_n367), .A3(KEYINPUT32), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n367), .B1(new_n358), .B2(KEYINPUT32), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n371), .B1(new_n477), .B2(new_n366), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n474), .B1(new_n478), .B2(new_n380), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n385), .A2(KEYINPUT74), .A3(new_n386), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n473), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n411), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n405), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(new_n406), .B2(new_n408), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n468), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n451), .A3(new_n450), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT84), .B(KEYINPUT35), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n481), .A2(new_n487), .A3(new_n276), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n399), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n404), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n399), .A2(KEYINPUT37), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n395), .A2(new_n398), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n405), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n495), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n494), .B1(new_n395), .B2(new_n398), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n404), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT38), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n486), .A2(new_n498), .A3(new_n469), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n422), .A2(new_n436), .A3(new_n438), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n440), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n448), .A2(new_n439), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT39), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n508), .A3(new_n440), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n417), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n507), .A2(KEYINPUT40), .A3(new_n417), .A4(new_n509), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n484), .A3(new_n513), .A4(new_n485), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n514), .A3(new_n276), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n272), .A2(new_n275), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n471), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n387), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n473), .A2(new_n518), .A3(new_n479), .A4(new_n480), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n515), .A2(new_n517), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n490), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G22gat), .Z(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n523), .A2(KEYINPUT88), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n523), .B2(KEYINPUT88), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n525), .B(new_n526), .C1(KEYINPUT16), .C2(new_n523), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(G8gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(G8gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT14), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT87), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT86), .B(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n533), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n540), .B(new_n544), .C1(KEYINPUT15), .C2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n543), .B2(new_n538), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n532), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n532), .B(new_n549), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n531), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n530), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n554), .B(new_n530), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n556), .B(KEYINPUT13), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n555), .A4(new_n556), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT85), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT11), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(new_n310), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT12), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n565), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G230gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n208), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(KEYINPUT9), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT89), .B(G57gat), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G64gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n401), .A2(G57gat), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G57gat), .B(G64gat), .Z(new_n583));
  AOI211_X1 g382(.A(new_n576), .B(new_n577), .C1(new_n583), .C2(KEYINPUT9), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT92), .A2(G85gat), .A3(G92gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n586), .A2(new_n587), .B1(new_n588), .B2(KEYINPUT8), .ZN(new_n589));
  OAI221_X1 g388(.A(new_n589), .B1(new_n587), .B2(new_n586), .C1(G85gat), .C2(G92gat), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n585), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n590), .B(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT94), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(KEYINPUT94), .A3(new_n585), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT10), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n585), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n575), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n598), .A2(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n574), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n309), .ZN(new_n608));
  INV_X1    g407(.A(G204gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT96), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n606), .A2(KEYINPUT95), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n606), .B2(KEYINPUT95), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n572), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n530), .B1(KEYINPUT21), .B2(new_n585), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n585), .A2(KEYINPUT21), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G127gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT90), .B(G155gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n624), .B(new_n627), .Z(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT91), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G162gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n596), .B1(new_n550), .B2(new_n552), .ZN(new_n633));
  NAND3_X1  g432(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(G190gat), .B(G218gat), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n554), .A2(new_n593), .B1(KEYINPUT93), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G134gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n636), .A2(KEYINPUT93), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G134gat), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n633), .A2(new_n642), .A3(new_n634), .A4(new_n637), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n641), .B1(new_n639), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n632), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n631), .A3(new_n644), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n628), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n522), .A2(new_n616), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n486), .A2(new_n469), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT97), .B(G1gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1324gat));
  AND2_X1   g456(.A1(new_n652), .A2(new_n484), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT16), .ZN(new_n659));
  INV_X1    g458(.A(G8gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n658), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT42), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(KEYINPUT42), .B2(new_n662), .ZN(G1325gat));
  AOI21_X1  g464(.A(G15gat), .B1(new_n652), .B2(new_n481), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n520), .B1(new_n518), .B2(new_n387), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT98), .Z(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n652), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n516), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT99), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT43), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(G22gat), .Z(G1327gat));
  AOI21_X1  g473(.A(new_n276), .B1(new_n653), .B2(new_n412), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n676), .A2(new_n515), .B1(new_n472), .B2(new_n489), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n616), .A2(new_n628), .ZN(new_n678));
  INV_X1    g477(.A(new_n650), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n533), .A3(new_n654), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT45), .Z(new_n682));
  INV_X1    g481(.A(new_n678), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n522), .B2(new_n650), .ZN(new_n685));
  AOI211_X1 g484(.A(KEYINPUT44), .B(new_n679), .C1(new_n490), .C2(new_n521), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT44), .B1(new_n677), .B2(new_n679), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n522), .A2(new_n684), .A3(new_n650), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n683), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n694), .A2(KEYINPUT101), .A3(new_n654), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT101), .B1(new_n694), .B2(new_n654), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n682), .B1(new_n697), .B2(G29gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT102), .ZN(G1328gat));
  AOI21_X1  g498(.A(new_n542), .B1(new_n694), .B2(new_n484), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n680), .A2(new_n542), .A3(new_n484), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n700), .A2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n680), .A2(new_n704), .A3(new_n481), .ZN(new_n705));
  INV_X1    g504(.A(new_n667), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT104), .Z(new_n708));
  OAI211_X1 g507(.A(KEYINPUT47), .B(new_n705), .C1(new_n708), .C2(new_n704), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n704), .B1(new_n694), .B2(new_n668), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n705), .B(KEYINPUT103), .Z(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n276), .B1(new_n688), .B2(new_n693), .ZN(new_n715));
  INV_X1    g514(.A(G50gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n692), .B1(new_n691), .B2(new_n683), .ZN(new_n718));
  AOI211_X1 g517(.A(KEYINPUT100), .B(new_n678), .C1(new_n689), .C2(new_n690), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n516), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n680), .A2(new_n716), .A3(new_n516), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n724), .ZN(new_n728));
  OAI21_X1  g527(.A(G50gat), .B1(new_n687), .B2(new_n276), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n722), .A3(KEYINPUT48), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT107), .Z(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n727), .A2(new_n734), .A3(new_n728), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1331gat));
  AND3_X1   g535(.A1(new_n522), .A2(new_n572), .A3(new_n651), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n614), .A2(new_n653), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n579), .B(KEYINPUT109), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n615), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n412), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT110), .Z(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n746), .B(new_n747), .Z(G1333gat));
  NAND3_X1  g547(.A1(new_n743), .A2(G71gat), .A3(new_n668), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT111), .Z(new_n750));
  XOR2_X1   g549(.A(new_n481), .B(KEYINPUT112), .Z(new_n751));
  AOI21_X1  g550(.A(G71gat), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g553(.A1(new_n614), .A2(new_n276), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  INV_X1    g556(.A(new_n628), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n565), .B(new_n570), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n522), .A3(new_n650), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT51), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT113), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n738), .A2(new_n416), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n691), .A2(new_n760), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n738), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n767), .A2(new_n768), .B1(new_n770), .B2(new_n416), .ZN(G1336gat));
  AND2_X1   g570(.A1(new_n769), .A2(new_n615), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n403), .B1(new_n772), .B2(new_n484), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n614), .A2(new_n412), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n403), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n762), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT52), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n767), .A2(new_n775), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(G1337gat));
  NAND2_X1  g579(.A1(new_n772), .A2(new_n668), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT114), .Z(new_n782));
  INV_X1    g581(.A(G99gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n615), .A2(new_n783), .A3(new_n481), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n782), .A2(new_n783), .B1(new_n767), .B2(new_n784), .ZN(G1338gat));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n755), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n516), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT115), .Z(new_n790));
  OAI221_X1 g589(.A(new_n786), .B1(new_n767), .B2(new_n788), .C1(new_n790), .C2(new_n787), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n762), .A2(new_n788), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(G106gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n786), .B2(new_n793), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n559), .A2(new_n562), .A3(new_n563), .A4(new_n570), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n560), .A2(new_n561), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n556), .B1(new_n553), .B2(new_n555), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n569), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n615), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n574), .B(new_n601), .C1(new_n604), .C2(KEYINPUT10), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n603), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n610), .B1(new_n603), .B2(KEYINPUT54), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n606), .A2(new_n610), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n603), .A2(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n603), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT55), .A4(new_n610), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n572), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n679), .ZN(new_n813));
  INV_X1    g612(.A(new_n811), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n650), .A2(new_n814), .A3(new_n800), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n758), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NOR4_X1   g615(.A1(new_n628), .A2(new_n759), .A3(new_n650), .A4(new_n615), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n795), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n817), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n650), .A2(new_n814), .A3(new_n800), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n679), .B2(new_n812), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n819), .B(KEYINPUT116), .C1(new_n821), .C2(new_n758), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n388), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n654), .A3(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n826), .A2(new_n412), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n572), .A2(new_n290), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT118), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n653), .A2(new_n484), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n276), .A3(new_n481), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n572), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(G1340gat));
  NAND3_X1  g635(.A1(new_n828), .A2(new_n280), .A3(new_n615), .ZN(new_n837));
  OAI21_X1  g636(.A(G120gat), .B1(new_n834), .B2(new_n614), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n834), .A2(new_n840), .A3(new_n628), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n828), .A2(new_n758), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n840), .ZN(G1342gat));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n642), .A3(new_n412), .A4(new_n827), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT56), .B1(new_n844), .B2(new_n679), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n846));
  OR3_X1    g645(.A1(new_n844), .A2(KEYINPUT56), .A3(new_n679), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(KEYINPUT56), .C1(new_n844), .C2(new_n679), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n834), .B2(new_n679), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n846), .A2(new_n847), .A3(new_n849), .A4(new_n850), .ZN(G1343gat));
  NAND2_X1  g650(.A1(new_n811), .A2(KEYINPUT121), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n806), .A2(new_n853), .A3(new_n807), .A4(new_n810), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n759), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n650), .B1(new_n855), .B2(new_n801), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n628), .B1(new_n856), .B2(new_n820), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT122), .B(new_n628), .C1(new_n856), .C2(new_n820), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n819), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n516), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n818), .A2(new_n822), .A3(new_n864), .A4(new_n516), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n706), .A2(new_n832), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT120), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n572), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n668), .A2(new_n276), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n833), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n759), .A2(new_n219), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT58), .ZN(G1344gat));
  AOI21_X1  g674(.A(new_n864), .B1(new_n861), .B2(new_n516), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n865), .A2(new_n867), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n614), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n221), .A2(new_n222), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(KEYINPUT59), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT123), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(new_n881), .C1(new_n869), .C2(new_n614), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n818), .A2(new_n516), .A3(new_n822), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n857), .A2(new_n819), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n864), .A3(new_n516), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n887), .A2(new_n615), .A3(new_n867), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G148gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT59), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n883), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n872), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n880), .A3(new_n615), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT124), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n893), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n869), .B2(new_n628), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n758), .A2(new_n233), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n872), .B2(new_n902), .ZN(G1346gat));
  AND2_X1   g702(.A1(new_n211), .A2(new_n213), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n905), .A3(new_n650), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n869), .A2(new_n679), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT125), .Z(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(new_n905), .ZN(G1347gat));
  NAND2_X1  g708(.A1(new_n823), .A2(new_n653), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n412), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n276), .A3(new_n751), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n572), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n823), .A2(new_n824), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n654), .A2(new_n412), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n759), .B1(new_n311), .B2(new_n312), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  OAI21_X1  g717(.A(G176gat), .B1(new_n912), .B2(new_n614), .ZN(new_n919));
  INV_X1    g718(.A(new_n910), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n920), .A2(new_n309), .A3(new_n824), .A4(new_n774), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n912), .B2(new_n628), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n758), .B1(new_n317), .B2(new_n316), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g725(.A1(new_n912), .A2(new_n679), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n927), .B2(new_n315), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(G190gat), .C1(new_n912), .C2(new_n679), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n914), .A2(new_n315), .A3(new_n650), .A4(new_n915), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT126), .B(new_n933), .C1(new_n927), .C2(new_n315), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n887), .A2(new_n889), .ZN(new_n936));
  INV_X1    g735(.A(new_n668), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n915), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n572), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n911), .A2(new_n871), .ZN(new_n942));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n759), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(G1352gat));
  NAND4_X1  g744(.A1(new_n920), .A2(new_n609), .A3(new_n774), .A4(new_n871), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT62), .Z(new_n947));
  NOR3_X1   g746(.A1(new_n936), .A2(new_n614), .A3(new_n938), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n609), .B2(new_n948), .ZN(G1353gat));
  AOI21_X1  g748(.A(new_n246), .B1(new_n939), .B2(new_n758), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n951));
  AND2_X1   g750(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n942), .A2(new_n246), .A3(new_n758), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G1354gat));
  AOI21_X1  g755(.A(G218gat), .B1(new_n942), .B2(new_n650), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n679), .A2(new_n247), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n939), .B2(new_n958), .ZN(G1355gat));
endmodule


