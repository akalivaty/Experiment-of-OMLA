//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1389,
    new_n1390;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  NAND2_X1  g0040(.A1(G33), .A2(G41), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n241), .A2(G1), .A3(G13), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G77), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G222), .A2(G1698), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT66), .B(G223), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(G1698), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n249), .B1(new_n252), .B2(new_n247), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  AND2_X1   g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n242), .A2(new_n258), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G190), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(new_n267), .B(KEYINPUT70), .Z(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(G200), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n273), .A2(KEYINPUT67), .A3(new_n212), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT67), .B1(new_n273), .B2(new_n212), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n205), .A2(G20), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G50), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G50), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n206), .B1(new_n201), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n206), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n277), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n282), .B(new_n291), .C1(G50), .C2(new_n278), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n292), .A2(new_n293), .B1(G200), .B2(new_n265), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n268), .A2(new_n272), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n267), .B(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT10), .B(new_n271), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n292), .B1(new_n264), .B2(G169), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(KEYINPUT68), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n301), .A2(KEYINPUT68), .B1(new_n303), .B2(new_n264), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT3), .B(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n261), .A2(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n308), .C1(G223), .C2(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n242), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n260), .B1(new_n226), .B2(new_n262), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G179), .B2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n273), .A2(new_n212), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G58), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n322), .B2(new_n201), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n288), .A2(G159), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n307), .B2(G20), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n247), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n325), .B1(new_n330), .B2(G68), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n319), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT76), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT74), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n244), .A2(new_n246), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n243), .A2(KEYINPUT74), .A3(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n328), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT75), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n244), .A2(new_n246), .A3(new_n335), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT75), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n328), .A4(new_n337), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n327), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n325), .B1(new_n343), .B2(G68), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n334), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n327), .ZN(new_n346));
  INV_X1    g0146(.A(new_n338), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n347), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g0148(.A(G68), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n325), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT76), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n333), .B1(new_n345), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n285), .B1(new_n205), .B2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n280), .A2(new_n355), .B1(new_n279), .B2(new_n285), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n317), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT18), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT76), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n334), .B(KEYINPUT16), .C1(new_n349), .C2(new_n350), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n332), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n313), .A2(G190), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n313), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n356), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n317), .C1(new_n354), .C2(new_n357), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n345), .A2(new_n353), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n357), .B1(new_n372), .B2(new_n332), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n359), .A2(new_n369), .A3(new_n371), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  INV_X1    g0176(.A(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G226), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n247), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n307), .A2(KEYINPUT72), .A3(G226), .A4(new_n377), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n307), .A2(G232), .A3(G1698), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n262), .A2(KEYINPUT73), .ZN(new_n386));
  INV_X1    g0186(.A(G238), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n262), .B2(KEYINPUT73), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n386), .A2(new_n388), .B1(new_n259), .B2(new_n257), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n385), .B2(new_n389), .ZN(new_n393));
  OAI21_X1  g0193(.A(G169), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n385), .A2(new_n389), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n391), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT14), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(G169), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(G179), .A3(new_n391), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n321), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n248), .B2(new_n286), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n277), .A2(KEYINPUT11), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n279), .A2(new_n321), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT12), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n279), .A2(new_n318), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(G68), .A3(new_n281), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT11), .B1(new_n277), .B2(new_n404), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n398), .A2(G200), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n397), .A2(G190), .A3(new_n391), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G244), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n260), .B1(new_n419), .B2(new_n262), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n307), .A2(G238), .A3(G1698), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n307), .A2(G232), .A3(new_n377), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n307), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n420), .B1(new_n424), .B2(new_n384), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G169), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n408), .A2(G77), .A3(new_n281), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G77), .B2(new_n278), .ZN(new_n428));
  INV_X1    g0228(.A(new_n285), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n286), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n318), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n425), .A2(KEYINPUT69), .A3(new_n303), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT69), .B1(new_n425), .B2(new_n303), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n425), .A2(G190), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n434), .B(new_n439), .C1(new_n364), .C2(new_n425), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n306), .A2(new_n375), .A3(new_n418), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT5), .B(G41), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n257), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n242), .ZN(new_n450));
  INV_X1    g0250(.A(G264), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G250), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n377), .ZN(new_n454));
  INV_X1    g0254(.A(G257), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n244), .A2(new_n454), .A3(new_n246), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G294), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n242), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(G200), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n384), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G264), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n457), .A2(new_n458), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n384), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n462), .A2(new_n464), .A3(G190), .A4(new_n446), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n244), .A2(new_n246), .A3(new_n206), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n307), .A2(new_n469), .A3(new_n206), .A4(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT81), .B(KEYINPUT24), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n206), .B2(G107), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n423), .A2(KEYINPUT23), .A3(G20), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n245), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n206), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n471), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n318), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n205), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n276), .A2(new_n278), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n423), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n279), .A2(new_n423), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT25), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n466), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT83), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT83), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n466), .A2(new_n481), .A3(new_n490), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n481), .A2(new_n487), .ZN(new_n492));
  OAI21_X1  g0292(.A(G169), .B1(new_n452), .B2(new_n459), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n462), .A2(new_n464), .A3(G179), .A4(new_n446), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n493), .B2(new_n494), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n489), .A2(new_n491), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n279), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n483), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g0302(.A(G107), .B1(new_n346), .B2(new_n348), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n504), .A2(new_n500), .A3(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(G97), .B(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n507), .A2(new_n206), .B1(new_n248), .B2(new_n289), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n502), .B1(new_n510), .B2(new_n318), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT78), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n419), .A2(G1698), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n244), .A3(new_n246), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT77), .A2(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n307), .A2(G250), .A3(G1698), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  INV_X1    g0318(.A(new_n515), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n513), .A3(new_n244), .A4(new_n246), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n384), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n449), .A2(G257), .A3(new_n242), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n446), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n512), .B1(new_n525), .B2(new_n266), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n449), .A2(new_n384), .A3(new_n255), .ZN(new_n527));
  AOI211_X1 g0327(.A(new_n527), .B(new_n523), .C1(new_n521), .C2(new_n384), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(KEYINPUT78), .A3(G190), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(G200), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n511), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n502), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n508), .B1(new_n343), .B2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n319), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n522), .A2(new_n303), .A3(new_n446), .A4(new_n524), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n314), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G257), .A2(G1698), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n377), .A2(G264), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n307), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT80), .B(G303), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n247), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n543), .A3(new_n384), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n449), .A2(G270), .A3(new_n242), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n446), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n319), .A2(new_n278), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n482), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n205), .A2(G13), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n476), .A2(G20), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n548), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n518), .B(new_n206), .C1(G33), .C2(new_n500), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n318), .A3(new_n551), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n547), .B(new_n558), .C1(new_n266), .C2(new_n546), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n546), .A2(G169), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n556), .ZN(new_n563));
  INV_X1    g0363(.A(new_n552), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n565), .A2(KEYINPUT21), .A3(G169), .A4(new_n546), .ZN(new_n566));
  AND4_X1   g0366(.A1(G179), .A2(new_n544), .A3(new_n446), .A4(new_n545), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n559), .A2(new_n562), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n387), .A2(new_n377), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n419), .A2(G1698), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n244), .A2(new_n570), .A3(new_n246), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n477), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n384), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n453), .B1(new_n205), .B2(G45), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n257), .A2(new_n444), .B1(new_n242), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n303), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT79), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n242), .B1(new_n572), .B2(new_n573), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n242), .A2(G274), .A3(new_n444), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n242), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT79), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n303), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n431), .A2(new_n278), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n206), .B1(new_n382), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n500), .A3(new_n423), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n244), .A2(new_n246), .A3(new_n206), .A4(G68), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n588), .B1(new_n286), .B2(new_n500), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n587), .B1(new_n595), .B2(new_n318), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n276), .A2(new_n278), .A3(new_n431), .A4(new_n482), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n314), .B1(new_n580), .B2(new_n583), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n579), .A2(new_n586), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G238), .A2(G1698), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n419), .B2(G1698), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n477), .B1(new_n602), .B2(new_n307), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n577), .B(G190), .C1(new_n603), .C2(new_n242), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n276), .A2(G87), .A3(new_n278), .A4(new_n482), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n604), .A2(new_n596), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(G200), .B1(new_n580), .B2(new_n583), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n569), .A2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n442), .A2(new_n499), .A3(new_n538), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n305), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT17), .B1(new_n373), .B2(new_n366), .ZN(new_n613));
  NOR4_X1   g0413(.A1(new_n354), .A2(new_n368), .A3(new_n357), .A4(new_n365), .ZN(new_n614));
  INV_X1    g0414(.A(new_n417), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(new_n438), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n613), .B(new_n614), .C1(new_n616), .C2(new_n414), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n362), .A2(new_n356), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n370), .B1(new_n618), .B2(new_n317), .ZN(new_n619));
  INV_X1    g0419(.A(new_n371), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n612), .B1(new_n623), .B2(new_n300), .ZN(new_n624));
  INV_X1    g0424(.A(new_n442), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT84), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n581), .A2(new_n582), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n581), .B2(new_n582), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n575), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n314), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n596), .A2(new_n597), .B1(new_n584), .B2(new_n303), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(G200), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n631), .A2(new_n632), .B1(new_n606), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n535), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n523), .B1(new_n521), .B2(new_n384), .ZN(new_n636));
  AOI21_X1  g0436(.A(G169), .B1(new_n636), .B2(new_n446), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n634), .A2(new_n638), .A3(new_n639), .A4(new_n534), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n598), .A2(new_n578), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n583), .A2(KEYINPUT84), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n627), .ZN(new_n643));
  AOI21_X1  g0443(.A(G169), .B1(new_n643), .B2(new_n575), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n535), .B1(new_n528), .B2(G169), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n511), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n600), .A2(new_n608), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT86), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n537), .B2(new_n609), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT86), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n640), .A4(new_n646), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n489), .A2(new_n491), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n531), .A2(new_n537), .A3(new_n634), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n493), .A2(new_n494), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n492), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n562), .A2(new_n566), .A3(new_n568), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n481), .A2(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT85), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n652), .A2(new_n655), .B1(new_n659), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n624), .B1(new_n625), .B2(new_n669), .ZN(G369));
  OR3_X1    g0470(.A1(new_n550), .A2(KEYINPUT27), .A3(G20), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT27), .B1(new_n550), .B2(G20), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT87), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n671), .A2(KEYINPUT87), .A3(G213), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(KEYINPUT88), .B(G343), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT89), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT89), .ZN(new_n680));
  INV_X1    g0480(.A(new_n678), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n675), .A2(new_n680), .A3(new_n676), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n492), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n499), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n498), .A2(new_n492), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n683), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n558), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n665), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n569), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n660), .A2(new_n683), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n499), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n689), .A2(new_n666), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n209), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n591), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n215), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n652), .A2(new_n655), .ZN(new_n708));
  INV_X1    g0508(.A(new_n658), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n656), .A3(new_n667), .A4(new_n664), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n683), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT92), .B1(new_n669), .B2(new_n683), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n665), .B1(new_n492), .B2(new_n498), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n657), .A2(new_n717), .A3(new_n658), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n649), .A2(new_n650), .A3(new_n639), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n364), .B1(new_n643), .B2(new_n575), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n604), .A2(new_n596), .A3(new_n605), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n641), .A2(new_n644), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(new_n511), .A3(new_n648), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n719), .B(new_n646), .C1(new_n639), .C2(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n689), .C1(new_n718), .C2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n499), .A2(new_n538), .A3(new_n610), .A4(new_n689), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n452), .A2(new_n459), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n567), .A2(new_n727), .A3(new_n636), .A4(new_n584), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT90), .B1(new_n528), .B2(new_n727), .ZN(new_n731));
  INV_X1    g0531(.A(new_n727), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT90), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n525), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n630), .A2(new_n303), .A3(new_n546), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n728), .A2(new_n729), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n689), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n728), .A2(KEYINPUT91), .A3(new_n729), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT91), .B1(new_n728), .B2(new_n729), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n689), .B1(new_n745), .B2(new_n737), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n726), .B(new_n742), .C1(KEYINPUT31), .C2(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n716), .A2(new_n725), .B1(G330), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n707), .B1(new_n748), .B2(G1), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT93), .ZN(G364));
  INV_X1    g0550(.A(G13), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(new_n443), .A3(G20), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT94), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n702), .A2(new_n753), .A3(new_n205), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n209), .A2(new_n307), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n209), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n701), .A2(new_n307), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n215), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(new_n443), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n236), .A2(new_n443), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n757), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n212), .B1(G20), .B2(new_n314), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n754), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n206), .A2(G179), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n206), .A2(new_n303), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT95), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT95), .B1(new_n206), .B2(new_n303), .ZN(new_n781));
  AND3_X1   g0581(.A1(new_n780), .A2(new_n781), .A3(new_n772), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n777), .A2(G329), .B1(new_n782), .B2(G311), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n266), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n303), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n785), .A2(G326), .B1(new_n788), .B2(G294), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n778), .A2(new_n266), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(G303), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n771), .A2(new_n266), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n247), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n780), .A2(new_n786), .A3(new_n781), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(new_n800), .B2(G322), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n783), .A2(new_n789), .A3(new_n795), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n307), .B1(new_n790), .B2(new_n321), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(new_n423), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G87), .B2(new_n794), .ZN(new_n805));
  INV_X1    g0605(.A(new_n788), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n283), .B2(new_n784), .C1(new_n500), .C2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n803), .B(new_n807), .C1(G77), .C2(new_n782), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n799), .B(KEYINPUT96), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n320), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n777), .A2(G159), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT32), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n802), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n770), .B1(new_n813), .B2(new_n767), .ZN(new_n814));
  INV_X1    g0614(.A(new_n766), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n692), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n754), .B1(new_n692), .B2(G330), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G330), .B2(new_n692), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  AOI22_X1  g0620(.A1(new_n777), .A2(G311), .B1(new_n782), .B2(G116), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n247), .B1(new_n806), .B2(new_n500), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G294), .B2(new_n800), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n796), .A2(new_n590), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G107), .B2(new_n794), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n791), .A2(G283), .B1(new_n785), .B2(G303), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n821), .A2(new_n823), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n791), .A2(G150), .B1(new_n785), .B2(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  INV_X1    g0629(.A(new_n782), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n828), .B1(new_n829), .B2(new_n830), .C1(new_n809), .C2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT98), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n777), .A2(G132), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n247), .B1(new_n788), .B2(G58), .ZN(new_n836));
  INV_X1    g0636(.A(new_n796), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n794), .A2(G50), .B1(new_n837), .B2(G68), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n827), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n767), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n433), .A2(new_n318), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n683), .B1(new_n843), .B2(new_n428), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n438), .A2(new_n844), .A3(new_n440), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n438), .B2(new_n440), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n764), .ZN(new_n848));
  INV_X1    g0648(.A(new_n754), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n767), .A2(new_n764), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n248), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n842), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n713), .A2(new_n714), .A3(new_n847), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n645), .B1(new_n723), .B2(new_n639), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n654), .B1(new_n854), .B2(new_n653), .ZN(new_n855));
  INV_X1    g0655(.A(new_n655), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n710), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n441), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n689), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n747), .A2(G330), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT99), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n861), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n862), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n864), .B2(new_n866), .ZN(G384));
  AOI21_X1  g0667(.A(new_n205), .B1(G13), .B2(new_n206), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n413), .A2(new_n683), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n414), .A2(new_n417), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n413), .B(new_n683), .C1(new_n615), .C2(new_n402), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n847), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n745), .A2(new_n737), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n683), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n740), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n746), .A2(KEYINPUT31), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n726), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n872), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(new_n677), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n354), .B2(new_n357), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n358), .A2(new_n882), .A3(new_n367), .A4(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n354), .A2(new_n357), .A3(new_n365), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n276), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(KEYINPUT16), .B2(new_n331), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n316), .A2(new_n677), .B1(new_n887), .B2(new_n356), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n356), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n881), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI221_X4 g0692(.A(new_n880), .B1(new_n884), .B2(new_n889), .C1(new_n375), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n375), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n884), .A2(new_n889), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n879), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n872), .A2(new_n877), .ZN(new_n898));
  INV_X1    g0698(.A(new_n882), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n375), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n358), .A2(new_n882), .A3(new_n367), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n884), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n880), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n898), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n897), .B1(new_n907), .B2(new_n878), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n442), .A3(new_n877), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n872), .A2(new_n877), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n900), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n893), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n613), .A2(new_n614), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n891), .B1(new_n621), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n895), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n880), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n906), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n912), .A2(KEYINPUT40), .B1(new_n917), .B2(new_n879), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n442), .A2(new_n877), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n909), .A2(G330), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT100), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n870), .A2(new_n871), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n438), .A2(new_n683), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n859), .B2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n928), .A2(new_n917), .B1(new_n622), .B2(new_n677), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n893), .B2(new_n911), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n402), .A2(new_n413), .A3(new_n689), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n716), .A2(new_n442), .A3(new_n725), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n624), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n868), .B1(new_n923), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n923), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(new_n507), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(KEYINPUT35), .ZN(new_n944));
  NOR4_X1   g0744(.A1(new_n943), .A2(new_n944), .A3(new_n214), .A4(new_n476), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  OR3_X1    g0746(.A1(new_n215), .A2(new_n248), .A3(new_n322), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n283), .A2(G68), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n751), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n946), .A3(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n796), .A2(new_n500), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G294), .B2(new_n791), .ZN(new_n953));
  INV_X1    g0753(.A(G311), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n784), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT46), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n793), .A2(new_n476), .B1(KEYINPUT107), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT107), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n809), .A2(new_n542), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n307), .B1(new_n788), .B2(G107), .ZN(new_n962));
  INV_X1    g0762(.A(G317), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n962), .B1(new_n776), .B2(new_n963), .C1(new_n797), .C2(new_n830), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n796), .A2(new_n248), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G68), .B2(new_n788), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n831), .B2(new_n784), .C1(new_n829), .C2(new_n790), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n307), .B1(new_n320), .B2(new_n793), .C1(new_n830), .C2(new_n283), .ZN(new_n969));
  INV_X1    g0769(.A(G137), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n776), .A2(new_n970), .B1(new_n799), .B2(new_n287), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT47), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n767), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n596), .A2(new_n605), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n683), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n634), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n646), .B2(new_n977), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(new_n815), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n768), .B1(new_n209), .B2(new_n432), .C1(new_n759), .C2(new_n232), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n982), .A2(new_n983), .A3(new_n849), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n975), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT102), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n683), .A2(new_n534), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n531), .A2(new_n537), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n649), .A2(new_n683), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n987), .B1(new_n992), .B2(new_n697), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(KEYINPUT42), .A3(new_n499), .A4(new_n696), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n498), .A2(new_n492), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n537), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n993), .A2(new_n994), .B1(new_n689), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT101), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(KEYINPUT101), .A3(new_n998), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT103), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n979), .B(KEYINPUT43), .Z(new_n1006));
  AND2_X1   g0806(.A1(new_n993), .A2(new_n994), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n996), .A2(new_n689), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1006), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT103), .B1(new_n997), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n986), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1014), .A2(new_n1003), .A3(KEYINPUT102), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1013), .A2(new_n1015), .B1(new_n695), .B2(new_n992), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1004), .A2(new_n986), .A3(new_n1012), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT102), .B1(new_n1014), .B2(new_n1003), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n695), .A2(new_n992), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n753), .A2(new_n205), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT104), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n992), .B1(new_n1024), .B2(KEYINPUT44), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(KEYINPUT44), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n1025), .A2(new_n699), .A3(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(KEYINPUT44), .C1(new_n699), .C2(new_n991), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n697), .A2(new_n698), .A3(new_n991), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT45), .ZN(new_n1031));
  OAI211_X1 g0831(.A(KEYINPUT105), .B(new_n694), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n694), .A2(KEYINPUT105), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n1028), .A4(new_n1027), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n697), .B1(new_n687), .B2(new_n696), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(new_n693), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n748), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n702), .B(KEYINPUT41), .Z(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1023), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n985), .B1(new_n1021), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(KEYINPUT108), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT108), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1045), .B(new_n985), .C1(new_n1021), .C2(new_n1042), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1046), .ZN(G387));
  NAND2_X1  g0847(.A1(new_n716), .A2(new_n725), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n861), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n1038), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1038), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n748), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n702), .A3(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n755), .A2(new_n704), .B1(G107), .B2(new_n209), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n229), .A2(G45), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT109), .Z(new_n1056));
  NOR3_X1   g0856(.A1(new_n285), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT50), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n429), .B2(new_n283), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n704), .B(new_n443), .C1(new_n321), .C2(new_n248), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1057), .B(new_n1059), .C1(new_n1061), .C2(KEYINPUT110), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(KEYINPUT110), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n759), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1054), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n247), .B(new_n952), .C1(new_n782), .C2(G68), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n283), .B2(new_n799), .C1(new_n287), .C2(new_n776), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n806), .A2(new_n432), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n784), .A2(new_n829), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n794), .A2(G77), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n285), .B2(new_n790), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n777), .A2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n247), .B1(new_n796), .B2(new_n476), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n791), .A2(G311), .B1(new_n785), .B2(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n542), .B2(new_n830), .C1(new_n809), .C2(new_n963), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  INV_X1    g0879(.A(G294), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n806), .A2(new_n797), .B1(new_n793), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1073), .B(new_n1074), .C1(new_n1082), .C2(KEYINPUT49), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1082), .A2(KEYINPUT49), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1072), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n767), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n754), .B1(new_n769), .B2(new_n1065), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n688), .B2(new_n766), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1051), .B2(new_n1023), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1053), .A2(new_n1089), .ZN(G393));
  NOR2_X1   g0890(.A1(new_n1052), .A2(new_n1036), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n703), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n694), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1033), .A2(new_n695), .A3(new_n1028), .A4(new_n1027), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1052), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(KEYINPUT111), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT111), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1052), .B2(new_n1095), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1093), .A2(new_n1023), .A3(new_n1094), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n768), .B1(new_n500), .B2(new_n209), .C1(new_n759), .C2(new_n239), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n754), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n793), .A2(new_n321), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n806), .A2(new_n248), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G50), .C2(new_n791), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n247), .B(new_n824), .C1(new_n782), .C2(new_n429), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n831), .C2(new_n776), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n799), .A2(new_n829), .B1(new_n287), .B2(new_n784), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT51), .Z(new_n1110));
  AOI211_X1 g0910(.A(new_n307), .B(new_n804), .C1(new_n777), .C2(G322), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n790), .A2(new_n542), .B1(new_n793), .B2(new_n797), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G116), .B2(new_n788), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n1080), .C2(new_n830), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n799), .A2(new_n954), .B1(new_n963), .B2(new_n784), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT52), .Z(new_n1116));
  OAI22_X1  g0916(.A1(new_n1108), .A2(new_n1110), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1103), .B1(new_n1117), .B2(new_n767), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n991), .B2(new_n815), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1101), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1100), .A2(new_n1121), .ZN(G390));
  NAND3_X1  g0922(.A1(new_n442), .A2(G330), .A3(new_n877), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n937), .A2(new_n624), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n847), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n742), .B1(new_n746), .B2(KEYINPUT31), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n726), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n1125), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n925), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n872), .A2(new_n877), .A3(G330), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1129), .A2(new_n1130), .B1(new_n859), .B2(new_n927), .ZN(new_n1131));
  AND4_X1   g0931(.A1(G330), .A2(new_n747), .A3(new_n924), .A4(new_n1125), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n877), .A2(G330), .A3(new_n1125), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n925), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n858), .B(new_n689), .C1(new_n718), .C2(new_n724), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT112), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n927), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1135), .B2(new_n927), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1131), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT113), .B1(new_n928), .B2(new_n934), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n931), .A2(new_n932), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT113), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n926), .B1(new_n711), .B2(new_n858), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n933), .C1(new_n1146), .C2(new_n925), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1137), .A2(new_n1138), .A3(new_n925), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n933), .B1(new_n893), .B2(new_n911), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1132), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1130), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1142), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n933), .B1(new_n1146), .B2(new_n925), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(KEYINPUT113), .B1(new_n931), .B2(new_n932), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1159), .B2(new_n1147), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1156), .B(new_n1141), .C1(new_n1160), .C2(new_n1130), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n702), .A3(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1156), .B(new_n1023), .C1(new_n1160), .C2(new_n1130), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1144), .A2(new_n764), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n776), .A2(new_n1080), .B1(new_n321), .B2(new_n796), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT114), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n785), .A2(G283), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1105), .B1(G107), .B2(new_n791), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n247), .B1(new_n590), .B2(new_n793), .C1(new_n799), .C2(new_n476), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G97), .B2(new_n782), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  INV_X1    g0972(.A(G132), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n830), .A2(new_n1172), .B1(new_n1173), .B2(new_n799), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n806), .A2(new_n829), .B1(new_n790), .B2(new_n970), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G128), .B2(new_n785), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n307), .B1(new_n796), .B2(new_n283), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n777), .B2(G125), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n793), .A2(new_n287), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT53), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1175), .A2(new_n1177), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1086), .B1(new_n1171), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n849), .B(new_n1183), .C1(new_n285), .C2(new_n850), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1164), .A2(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1163), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT115), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1162), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1162), .B2(new_n1186), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(G378));
  NAND2_X1  g0990(.A1(new_n292), .A2(new_n881), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT118), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n612), .B1(new_n296), .B2(new_n299), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1193), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n306), .A2(new_n1195), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT119), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G330), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n918), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT119), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1202), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1192), .B1(new_n1201), .B2(new_n1197), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n908), .B2(G330), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n936), .B1(new_n1205), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1203), .B1(new_n918), .B2(new_n1204), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n936), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n908), .A2(G330), .A3(new_n1209), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n764), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n850), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n754), .B1(G50), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n307), .A2(G41), .ZN(new_n1220));
  INV_X1    g1020(.A(G41), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G50), .B(new_n1220), .C1(new_n245), .C2(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n776), .A2(new_n797), .B1(new_n799), .B2(new_n423), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n431), .B2(new_n782), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1070), .A2(KEYINPUT116), .A3(new_n1220), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT116), .B1(new_n1070), .B2(new_n1220), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n806), .A2(new_n321), .B1(new_n784), .B2(new_n476), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n790), .A2(new_n500), .B1(new_n796), .B2(new_n320), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1224), .A2(new_n1225), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1222), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1172), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n785), .A2(G125), .B1(new_n794), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n287), .B2(new_n806), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n782), .A2(G137), .B1(G132), .B2(new_n791), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT117), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1235), .B(new_n1237), .C1(G128), .C2(new_n800), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n245), .B(new_n1221), .C1(new_n796), .C2(new_n829), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n777), .B2(G124), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT59), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1242), .B1(new_n1238), .B2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1232), .B1(new_n1231), .B2(new_n1230), .C1(new_n1240), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1219), .B1(new_n1245), .B2(new_n767), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1216), .A2(new_n1023), .B1(new_n1217), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1124), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1161), .A2(new_n1248), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1213), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n702), .B1(new_n1249), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1161), .A2(new_n1248), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1216), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1247), .B1(new_n1253), .B2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1142), .A2(new_n1041), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n849), .B1(new_n321), .B2(new_n850), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n806), .A2(new_n283), .B1(new_n793), .B2(new_n829), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n785), .A2(G132), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT120), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1260), .B(new_n1262), .C1(new_n791), .C2(new_n1233), .ZN(new_n1263));
  INV_X1    g1063(.A(G128), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n307), .B1(new_n320), .B2(new_n796), .C1(new_n776), .C2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G150), .B2(new_n782), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1263), .B(new_n1266), .C1(new_n970), .C2(new_n809), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n777), .A2(G303), .B1(new_n782), .B2(G107), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1068), .B1(G294), .B2(new_n785), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G116), .A2(new_n791), .B1(new_n794), .B2(G97), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n307), .B(new_n966), .C1(new_n800), .C2(G283), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT121), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n767), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1273), .A2(KEYINPUT121), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1259), .B1(new_n1275), .B2(new_n1276), .C1(new_n924), .C2(new_n765), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1140), .B2(new_n1022), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1258), .A2(new_n1279), .ZN(G381));
  XNOR2_X1  g1080(.A(new_n1096), .B(KEYINPUT111), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1120), .B1(new_n1281), .B2(new_n1092), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1285), .A2(G381), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1162), .A2(new_n1186), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G387), .A2(new_n1286), .A3(new_n1287), .A4(G375), .ZN(G407));
  NAND2_X1  g1088(.A1(new_n1216), .A2(new_n1023), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1217), .A2(new_n1246), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1254), .A2(new_n1216), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT57), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n703), .B1(new_n1295), .B2(new_n1254), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1291), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1287), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n678), .A2(G213), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT122), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G407), .A2(G213), .A3(new_n1301), .ZN(G409));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT124), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n985), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1020), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1019), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1042), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1305), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1310), .B2(G390), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1282), .A2(new_n1043), .A3(KEYINPUT124), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(G390), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(new_n819), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1044), .A2(new_n1046), .A3(new_n1282), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1315), .B1(new_n1310), .B2(G390), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT125), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1316), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1247), .B1(new_n1292), .B2(new_n1040), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1298), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1287), .A2(KEYINPUT115), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1162), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1325), .B1(new_n1328), .B2(G375), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1300), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1142), .A2(new_n702), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT123), .B1(new_n1124), .B2(new_n1140), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1332), .A2(KEYINPUT60), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(KEYINPUT60), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1331), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1336), .A2(new_n1283), .A3(new_n1278), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1332), .A2(KEYINPUT60), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n702), .B(new_n1142), .C1(new_n1338), .C2(new_n1333), .ZN(new_n1339));
  AOI21_X1  g1139(.A(G384), .B1(new_n1339), .B2(new_n1279), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1337), .A2(new_n1340), .ZN(new_n1341));
  AND4_X1   g1141(.A1(new_n1323), .A2(new_n1329), .A3(new_n1330), .A4(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1295), .A2(new_n1254), .ZN(new_n1343));
  AOI22_X1  g1143(.A1(new_n1161), .A2(new_n1248), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1343), .B(new_n702), .C1(KEYINPUT57), .C2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1345), .A2(new_n1326), .A3(new_n1327), .A4(new_n1247), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1300), .B1(new_n1346), .B2(new_n1325), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1323), .B1(new_n1347), .B2(new_n1341), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1342), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT61), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1300), .A2(G2897), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1283), .B1(new_n1336), .B2(new_n1278), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1339), .A2(G384), .A3(new_n1279), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1351), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1352), .A2(new_n1353), .A3(new_n1351), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1350), .B1(new_n1347), .B2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT126), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1322), .B1(new_n1349), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1351), .ZN(new_n1362));
  NOR3_X1   g1162(.A1(new_n1337), .A2(new_n1340), .A3(new_n1362), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1363), .A2(new_n1354), .ZN(new_n1364));
  AOI22_X1  g1164(.A1(G378), .A2(new_n1297), .B1(new_n1298), .B2(new_n1324), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1364), .B1(new_n1365), .B2(new_n1300), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1316), .B(new_n1359), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1366), .A2(new_n1367), .A3(new_n1350), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1329), .A2(new_n1330), .A3(new_n1341), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT63), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1347), .A2(KEYINPUT63), .A3(new_n1341), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1368), .B1(new_n1373), .B2(new_n1322), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1303), .B1(new_n1361), .B2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1372), .ZN(new_n1376));
  AOI21_X1  g1176(.A(KEYINPUT63), .B1(new_n1347), .B2(new_n1341), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1322), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1378));
  INV_X1    g1178(.A(new_n1368), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(new_n1322), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1369), .A2(KEYINPUT62), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1347), .A2(new_n1323), .A3(new_n1341), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1184(.A(KEYINPUT126), .B1(new_n1366), .B2(new_n1350), .ZN(new_n1385));
  OAI21_X1  g1185(.A(new_n1381), .B1(new_n1384), .B2(new_n1385), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1380), .A2(new_n1386), .A3(KEYINPUT127), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1375), .A2(new_n1387), .ZN(G405));
  OAI21_X1  g1188(.A(new_n1346), .B1(new_n1287), .B2(new_n1297), .ZN(new_n1389));
  XNOR2_X1  g1189(.A(new_n1389), .B(new_n1341), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(new_n1390), .B(new_n1381), .ZN(G402));
endmodule


