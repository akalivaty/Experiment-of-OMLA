//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT69), .Z(G261));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR3_X1   g035(.A1(new_n456), .A2(KEYINPUT70), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n455), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G2106), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT70), .B1(new_n456), .B2(new_n460), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n473), .A2(new_n475), .A3(G137), .A4(new_n467), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n475), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(KEYINPUT71), .A3(G136), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n468), .A2(new_n467), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n480), .A2(new_n467), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n482), .A2(new_n486), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n503), .A2(new_n468), .A3(G138), .A4(new_n467), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n467), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n500), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n498), .B1(new_n504), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n513), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n522), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n512), .A2(new_n517), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n509), .A2(new_n511), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n509), .B2(new_n511), .ZN(new_n534));
  OAI211_X1 g109(.A(G63), .B(G651), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT74), .B(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n517), .A2(G543), .A3(new_n537), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n536), .B1(new_n535), .B2(new_n538), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n528), .B(new_n531), .C1(new_n539), .C2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n518), .A2(new_n543), .B1(new_n520), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n509), .A2(new_n511), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT73), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n509), .A2(new_n511), .A3(new_n532), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G64), .ZN(new_n550));
  INV_X1    g125(.A(G77), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n551), .B2(new_n508), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n545), .B1(new_n552), .B2(G651), .ZN(G171));
  INV_X1    g128(.A(new_n520), .ZN(new_n554));
  AOI22_X1  g129(.A1(G43), .A2(new_n554), .B1(new_n529), .B2(G81), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n549), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n513), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n555), .B(new_n559), .C1(new_n513), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n518), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n512), .A2(new_n517), .A3(KEYINPUT78), .A4(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n520), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n517), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n513), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n572), .A2(new_n577), .A3(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  OAI21_X1  g156(.A(G651), .B1(new_n549), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n529), .A2(G87), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n514), .A2(new_n516), .A3(G49), .A4(G543), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(G288));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n518), .A2(new_n588), .B1(new_n520), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n513), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n549), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n513), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n518), .A2(new_n598), .B1(new_n520), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n529), .A2(KEYINPUT81), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n518), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n606), .B1(new_n605), .B2(new_n609), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n615));
  INV_X1    g190(.A(G79), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n616), .A2(new_n508), .A3(KEYINPUT82), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(new_n616), .B2(new_n508), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n546), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n554), .A2(G54), .B1(new_n620), .B2(G651), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n613), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n603), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n603), .B1(new_n622), .B2(G868), .ZN(G321));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G299), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G168), .B2(new_n625), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(G168), .B2(new_n625), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n487), .A2(G123), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n481), .A2(G135), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n639));
  AND3_X1   g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(G156));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT15), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G2435), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT15), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(G2435), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n652), .A2(new_n656), .A3(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n657), .A2(new_n658), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n658), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1341), .B(G1348), .Z(new_n669));
  AOI21_X1  g244(.A(new_n648), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n671), .A3(new_n667), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g249(.A1(new_n664), .A2(KEYINPUT86), .A3(new_n671), .A4(new_n667), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n678));
  NAND4_X1  g253(.A1(new_n670), .A2(new_n674), .A3(new_n678), .A4(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n686), .B1(new_n690), .B2(KEYINPUT17), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(new_n685), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n690), .A2(KEYINPUT17), .A3(new_n686), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G2096), .B(G2100), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(G227));
  XOR2_X1   g273(.A(G1971), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n705), .A2(new_n706), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n708), .B(new_n709), .C1(new_n706), .C2(new_n705), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n712), .B(new_n716), .ZN(G229));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n487), .A2(G119), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G131), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n467), .A2(G107), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(G29), .ZN(new_n725));
  MUX2_X1   g300(.A(new_n719), .B(new_n725), .S(KEYINPUT93), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n726), .B(new_n727), .Z(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n601), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(G22), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G166), .B2(new_n729), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT96), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1971), .ZN(new_n737));
  MUX2_X1   g312(.A(G6), .B(G305), .S(G16), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT32), .B(G1981), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT94), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT95), .B1(G16), .B2(G23), .ZN(new_n742));
  OR3_X1    g317(.A1(KEYINPUT95), .A2(G16), .A3(G23), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n742), .B(new_n743), .C1(G288), .C2(new_n729), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT33), .B(G1976), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n737), .A2(KEYINPUT34), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT34), .B1(new_n737), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n733), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT97), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n487), .A2(G128), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n481), .A2(G140), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n467), .A2(G116), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT98), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n718), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n770), .A2(new_n718), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G160), .B2(new_n718), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n769), .B1(new_n756), .B2(G11), .C1(G2084), .C2(new_n773), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n757), .B(new_n774), .C1(G2084), .C2(new_n773), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT104), .B(KEYINPUT23), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n729), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n718), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n718), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT103), .B(G2078), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n775), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G35), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G162), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT29), .Z(new_n788));
  INV_X1    g363(.A(G2090), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n481), .A2(KEYINPUT99), .A3(G139), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT99), .B1(new_n481), .B2(G139), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n793), .B1(new_n467), .B2(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n790), .A2(new_n791), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n729), .A2(G5), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G171), .B2(new_n729), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT102), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G21), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G168), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT101), .B(G1966), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(G28), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(G28), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n811), .A2(new_n812), .A3(new_n718), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n800), .A2(new_n804), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G4), .A2(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n622), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1348), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n785), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n487), .A2(G129), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT100), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n821));
  NAND3_X1  g396(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT26), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G141), .B2(new_n481), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G32), .B(new_n825), .S(G29), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT27), .B(G1996), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n751), .A2(new_n752), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n750), .A2(new_n829), .A3(new_n754), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n755), .A2(new_n818), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G16), .A2(G19), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n561), .B2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1341), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n640), .A2(G29), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n831), .A2(new_n834), .A3(new_n836), .ZN(G311));
  OR3_X1    g412(.A1(new_n831), .A2(new_n834), .A3(new_n836), .ZN(G150));
  AOI22_X1  g413(.A1(new_n549), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT105), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  AOI22_X1  g416(.A1(G55), .A2(new_n554), .B1(new_n529), .B2(G93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n561), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n557), .A3(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n622), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n845), .B1(new_n852), .B2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT106), .Z(G145));
  XNOR2_X1  g429(.A(new_n491), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n640), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n825), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n797), .B(new_n762), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n504), .A2(new_n506), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n493), .A2(KEYINPUT107), .A3(new_n497), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT107), .B1(new_n493), .B2(new_n497), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n643), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n857), .B(new_n864), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n487), .A2(G130), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n467), .A2(G118), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n724), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n857), .B(new_n864), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n871), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT40), .Z(G395));
  AND2_X1   g453(.A1(new_n846), .A2(new_n847), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n631), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n622), .A2(G299), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n613), .A2(new_n615), .A3(new_n621), .ZN(new_n882));
  INV_X1    g457(.A(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n885), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(new_n880), .ZN(new_n890));
  INV_X1    g465(.A(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n601), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G303), .B(G305), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT42), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(G868), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT108), .B1(new_n843), .B2(new_n625), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n896), .A2(KEYINPUT108), .A3(G868), .A4(new_n897), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G295));
  AND2_X1   g477(.A1(new_n900), .A2(new_n901), .ZN(G331));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  XNOR2_X1  g479(.A(G301), .B(G286), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n879), .A2(KEYINPUT109), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n848), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n848), .B2(new_n907), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n888), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n885), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n848), .A2(new_n907), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n894), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n874), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n888), .B2(new_n911), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n894), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n904), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n919), .B2(new_n894), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n885), .A2(new_n887), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT41), .B1(new_n881), .B2(new_n884), .ZN(new_n924));
  INV_X1    g499(.A(new_n908), .ZN(new_n925));
  OAI22_X1  g500(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n914), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n906), .A2(new_n885), .A3(new_n910), .A4(new_n908), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n894), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n930), .B(new_n894), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n922), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n921), .B1(new_n932), .B2(new_n904), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT44), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n922), .B(new_n904), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n918), .B2(new_n920), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n862), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(KEYINPUT111), .B(G40), .Z(new_n945));
  NOR3_X1   g520(.A1(new_n471), .A2(new_n478), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n825), .B(G1996), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n762), .B(G2067), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n724), .A2(new_n727), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n762), .A2(G2067), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n949), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n949), .B2(G1996), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n948), .B1(new_n825), .B2(new_n951), .ZN(new_n959));
  INV_X1    g534(.A(G1996), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n948), .A2(KEYINPUT46), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  AND2_X1   g538(.A1(new_n724), .A2(new_n727), .ZN(new_n964));
  NOR4_X1   g539(.A1(new_n950), .A2(new_n964), .A3(new_n953), .A4(new_n951), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n965), .A2(new_n949), .ZN(new_n966));
  NOR2_X1   g541(.A1(G290), .A2(G1986), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n948), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT48), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n956), .B(new_n963), .C1(new_n966), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT124), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n862), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(G160), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(G2078), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n973), .A2(G40), .A3(new_n944), .A4(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G2078), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n943), .B1(G164), .B2(G1384), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n972), .A2(new_n977), .A3(new_n946), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n974), .ZN(new_n980));
  INV_X1    g555(.A(new_n498), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n859), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n946), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n862), .A2(new_n983), .A3(new_n941), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT112), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n862), .A2(new_n987), .A3(new_n983), .A4(new_n941), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n976), .B(new_n980), .C1(G1961), .C2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n971), .B1(new_n990), .B2(G171), .ZN(new_n991));
  NOR3_X1   g566(.A1(G164), .A2(new_n943), .A3(G1384), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n943), .A2(new_n942), .B1(new_n992), .B2(KEYINPUT118), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n982), .A2(KEYINPUT45), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n947), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n975), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n980), .C1(G1961), .C2(new_n989), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT54), .B1(new_n998), .B2(G171), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n986), .A2(new_n988), .ZN(new_n1000));
  INV_X1    g575(.A(new_n984), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1002), .A2(new_n1003), .B1(new_n974), .B2(new_n979), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(KEYINPUT124), .A3(G301), .A4(new_n976), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n991), .A2(new_n999), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(G301), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1007), .B(KEYINPUT54), .C1(G301), .C2(new_n990), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(G2084), .B(new_n984), .C1(new_n986), .C2(new_n988), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n807), .B1(new_n993), .B2(new_n996), .ZN(new_n1011));
  AND3_X1   g586(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT121), .B1(G286), .B2(G8), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n1010), .A2(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1015));
  INV_X1    g590(.A(KEYINPUT123), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G286), .A2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(KEYINPUT123), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  INV_X1    g599(.A(G2084), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1000), .A2(new_n1025), .A3(new_n1001), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n498), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n493), .A2(KEYINPUT107), .A3(new_n497), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n859), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n994), .A2(new_n995), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n946), .B1(new_n992), .B2(KEYINPUT118), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n808), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1024), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1014), .B(new_n1015), .C1(new_n1023), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(new_n1038), .C1(new_n1039), .C2(new_n1024), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT61), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n982), .A2(new_n983), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1043), .B(new_n946), .C1(new_n1031), .C2(new_n983), .ZN(new_n1044));
  INV_X1    g619(.A(G1956), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G299), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n572), .A2(new_n577), .A3(new_n579), .A4(KEYINPUT57), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT56), .B(G2072), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n972), .A2(new_n946), .A3(new_n978), .A4(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1046), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1042), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1050), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1046), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT61), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1348), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n946), .A2(new_n862), .A3(new_n941), .A4(new_n768), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n622), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1064), .B(KEYINPUT120), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n882), .B(new_n1068), .C1(G1348), .C2(new_n989), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1062), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1068), .B(new_n1062), .C1(new_n989), .C2(G1348), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n972), .A2(new_n960), .A3(new_n946), .A4(new_n978), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n946), .A2(new_n862), .A3(new_n941), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n561), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1076), .B2(new_n561), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1071), .A2(new_n882), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1061), .A2(new_n1070), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1053), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1009), .B(new_n1041), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G301), .B1(new_n1004), .B2(new_n997), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1036), .A2(KEYINPUT62), .A3(new_n1040), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT113), .B(G2090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n989), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n972), .A2(new_n946), .A3(new_n978), .ZN(new_n1094));
  INV_X1    g669(.A(G1971), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1024), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n1098));
  OAI221_X1 g673(.A(G8), .B1(new_n1098), .B2(KEYINPUT55), .C1(new_n522), .C2(new_n524), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(KEYINPUT55), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n1100), .B(KEYINPUT115), .Z(new_n1101));
  XNOR2_X1  g676(.A(new_n1099), .B(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1096), .B1(new_n1044), .B2(new_n1091), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1104), .B2(G8), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n582), .A2(G1976), .A3(new_n583), .A4(new_n586), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1073), .A2(G8), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(KEYINPUT116), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1024), .B1(new_n1031), .B2(new_n946), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(KEYINPUT116), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1976), .ZN(new_n1114));
  NAND3_X1  g689(.A1(G288), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n591), .A2(new_n594), .A3(new_n714), .ZN(new_n1118));
  OAI21_X1  g693(.A(G1981), .B1(new_n590), .B2(new_n593), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT49), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(KEYINPUT49), .A3(new_n1119), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1111), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1116), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1117), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1103), .B(new_n1106), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1090), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1035), .A2(G168), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1126), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1116), .A2(new_n1117), .A3(new_n1124), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1105), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1131), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(KEYINPUT119), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1116), .A2(new_n1124), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1103), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1124), .A2(new_n1114), .A3(new_n891), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1118), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1111), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(new_n1138), .A3(new_n1103), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT63), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1140), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1129), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1986), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n965), .B1(new_n1151), .B2(new_n601), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n948), .B1(new_n1152), .B2(new_n967), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT125), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1127), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1140), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT125), .B(new_n1153), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n970), .B1(new_n1154), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g734(.A1(G229), .A2(new_n465), .ZN(new_n1161));
  AOI211_X1 g735(.A(G227), .B(new_n1161), .C1(new_n677), .C2(new_n679), .ZN(new_n1162));
  AOI21_X1  g736(.A(new_n877), .B1(new_n1162), .B2(KEYINPUT126), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1164));
  INV_X1    g738(.A(G227), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n680), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1166), .B2(new_n1161), .ZN(new_n1167));
  AND3_X1   g741(.A1(new_n1163), .A2(new_n937), .A3(new_n1167), .ZN(G308));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n937), .A3(new_n1167), .ZN(G225));
endmodule


