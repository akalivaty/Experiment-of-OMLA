

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753;

  AND2_X1 U365 ( .A1(n548), .A2(n547), .ZN(n557) );
  AND2_X1 U366 ( .A1(n596), .A2(n595), .ZN(n597) );
  INV_X1 U367 ( .A(n605), .ZN(n701) );
  INV_X1 U368 ( .A(G953), .ZN(n731) );
  XNOR2_X1 U369 ( .A(n536), .B(n520), .ZN(n575) );
  XNOR2_X2 U370 ( .A(n489), .B(n411), .ZN(n426) );
  XNOR2_X2 U371 ( .A(n609), .B(n608), .ZN(n753) );
  NAND2_X1 U372 ( .A1(n571), .A2(n573), .ZN(n692) );
  AND2_X1 U373 ( .A1(n361), .A2(n546), .ZN(n547) );
  AND2_X1 U374 ( .A1(n386), .A2(n384), .ZN(n383) );
  XNOR2_X1 U375 ( .A(n519), .B(n396), .ZN(n395) );
  NAND2_X1 U376 ( .A1(n347), .A2(n393), .ZN(n607) );
  XNOR2_X1 U377 ( .A(n600), .B(KEYINPUT105), .ZN(n675) );
  XNOR2_X1 U378 ( .A(n651), .B(n650), .ZN(n652) );
  AND2_X1 U379 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U380 ( .A(n441), .B(n440), .ZN(n571) );
  NAND2_X1 U381 ( .A1(n370), .A2(n475), .ZN(n369) );
  XNOR2_X1 U382 ( .A(n486), .B(n375), .ZN(n742) );
  XNOR2_X1 U383 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n407) );
  BUF_X1 U384 ( .A(n663), .Z(n343) );
  OR2_X2 U385 ( .A1(n575), .A2(n692), .ZN(n382) );
  OR2_X1 U386 ( .A1(n641), .A2(n369), .ZN(n368) );
  BUF_X1 U387 ( .A(n732), .Z(n344) );
  NOR2_X2 U388 ( .A1(n382), .A2(n535), .ZN(n381) );
  NAND2_X1 U389 ( .A1(n395), .A2(n535), .ZN(n528) );
  NOR2_X2 U390 ( .A1(n607), .A2(n586), .ZN(n673) );
  XNOR2_X2 U391 ( .A(n744), .B(n409), .ZN(n489) );
  XNOR2_X1 U392 ( .A(n353), .B(n435), .ZN(n635) );
  XNOR2_X1 U393 ( .A(n345), .B(n434), .ZN(n435) );
  XNOR2_X1 U394 ( .A(n436), .B(n742), .ZN(n353) );
  XNOR2_X1 U395 ( .A(n461), .B(n374), .ZN(n656) );
  XNOR2_X1 U396 ( .A(n376), .B(n742), .ZN(n374) );
  INV_X1 U397 ( .A(KEYINPUT22), .ZN(n396) );
  INV_X1 U398 ( .A(KEYINPUT6), .ZN(n520) );
  INV_X1 U399 ( .A(n666), .ZN(n363) );
  XNOR2_X1 U400 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n428) );
  XNOR2_X1 U401 ( .A(G119), .B(G128), .ZN(n430) );
  XNOR2_X1 U402 ( .A(n454), .B(n377), .ZN(n376) );
  XNOR2_X1 U403 ( .A(n455), .B(n453), .ZN(n377) );
  XNOR2_X1 U404 ( .A(G140), .B(KEYINPUT10), .ZN(n375) );
  XNOR2_X1 U405 ( .A(G110), .B(G104), .ZN(n480) );
  XNOR2_X1 U406 ( .A(n381), .B(n549), .ZN(n387) );
  OR2_X1 U407 ( .A1(n627), .A2(G902), .ZN(n427) );
  NOR2_X1 U408 ( .A1(n623), .A2(n401), .ZN(n400) );
  AND2_X1 U409 ( .A1(n621), .A2(n402), .ZN(n401) );
  XNOR2_X1 U410 ( .A(n378), .B(KEYINPUT107), .ZN(n576) );
  NAND2_X1 U411 ( .A1(n379), .A2(n675), .ZN(n378) );
  NAND2_X1 U412 ( .A1(n383), .A2(n390), .ZN(n553) );
  XNOR2_X1 U413 ( .A(n463), .B(n462), .ZN(n543) );
  XNOR2_X1 U414 ( .A(n642), .B(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U415 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U416 ( .A(n656), .B(KEYINPUT59), .ZN(n657) );
  XNOR2_X1 U417 ( .A(n627), .B(n626), .ZN(n628) );
  AND2_X1 U418 ( .A1(n630), .A2(G953), .ZN(n726) );
  NAND2_X1 U419 ( .A1(n360), .A2(n523), .ZN(n546) );
  INV_X1 U420 ( .A(n528), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n720) );
  INV_X1 U422 ( .A(KEYINPUT119), .ZN(n354) );
  XOR2_X1 U423 ( .A(n431), .B(n430), .Z(n345) );
  NOR2_X1 U424 ( .A1(n543), .A2(n514), .ZN(n346) );
  XOR2_X1 U425 ( .A(n583), .B(n582), .Z(n347) );
  AND2_X1 U426 ( .A1(n525), .A2(n575), .ZN(n348) );
  XOR2_X1 U427 ( .A(n503), .B(KEYINPUT19), .Z(n349) );
  NOR2_X1 U428 ( .A1(n402), .A2(n621), .ZN(n350) );
  INV_X1 U429 ( .A(KEYINPUT80), .ZN(n402) );
  NAND2_X1 U430 ( .A1(n732), .A2(n745), .ZN(n351) );
  AND2_X2 U431 ( .A1(n620), .A2(n619), .ZN(n745) );
  NAND2_X1 U432 ( .A1(n357), .A2(KEYINPUT2), .ZN(n356) );
  NOR2_X1 U433 ( .A1(n703), .A2(n686), .ZN(n517) );
  NAND2_X2 U434 ( .A1(n352), .A2(n359), .ZN(n358) );
  AND2_X2 U435 ( .A1(n397), .A2(n400), .ZN(n352) );
  INV_X1 U436 ( .A(n351), .ZN(n357) );
  XNOR2_X2 U437 ( .A(n413), .B(n412), .ZN(n478) );
  AND2_X1 U438 ( .A1(n745), .A2(n350), .ZN(n399) );
  INV_X1 U439 ( .A(n692), .ZN(n391) );
  NAND2_X1 U440 ( .A1(n719), .A2(n718), .ZN(n355) );
  AND2_X4 U441 ( .A1(n358), .A2(n356), .ZN(n722) );
  INV_X1 U442 ( .A(n398), .ZN(n359) );
  NAND2_X1 U443 ( .A1(n732), .A2(n745), .ZN(n624) );
  AND2_X1 U444 ( .A1(n732), .A2(n399), .ZN(n398) );
  XNOR2_X2 U445 ( .A(n365), .B(n568), .ZN(n732) );
  NAND2_X1 U446 ( .A1(n362), .A2(n545), .ZN(n361) );
  NAND2_X1 U447 ( .A1(n364), .A2(n363), .ZN(n362) );
  INV_X1 U448 ( .A(n678), .ZN(n364) );
  XNOR2_X2 U449 ( .A(n538), .B(KEYINPUT31), .ZN(n678) );
  NAND2_X1 U450 ( .A1(n366), .A2(n567), .ZN(n365) );
  XNOR2_X1 U451 ( .A(n367), .B(n558), .ZN(n366) );
  NAND2_X1 U452 ( .A1(n556), .A2(n557), .ZN(n367) );
  NAND2_X4 U453 ( .A1(n371), .A2(n368), .ZN(n536) );
  INV_X1 U454 ( .A(n418), .ZN(n370) );
  NAND2_X1 U455 ( .A1(n418), .A2(G902), .ZN(n372) );
  NAND2_X1 U456 ( .A1(n641), .A2(n418), .ZN(n373) );
  XNOR2_X2 U457 ( .A(n513), .B(n512), .ZN(n534) );
  AND2_X1 U458 ( .A1(n380), .A2(n580), .ZN(n379) );
  INV_X1 U459 ( .A(n575), .ZN(n380) );
  INV_X1 U460 ( .A(n535), .ZN(n578) );
  INV_X1 U461 ( .A(n387), .ZN(n709) );
  AND2_X1 U462 ( .A1(n385), .A2(n346), .ZN(n384) );
  NAND2_X1 U463 ( .A1(n550), .A2(KEYINPUT34), .ZN(n385) );
  NAND2_X1 U464 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U465 ( .A1(n550), .A2(KEYINPUT34), .ZN(n388) );
  XNOR2_X2 U466 ( .A(n389), .B(G143), .ZN(n472) );
  XNOR2_X2 U467 ( .A(G128), .B(KEYINPUT66), .ZN(n389) );
  NAND2_X1 U468 ( .A1(n709), .A2(KEYINPUT34), .ZN(n390) );
  NAND2_X1 U469 ( .A1(n393), .A2(n391), .ZN(n539) );
  XNOR2_X2 U470 ( .A(n393), .B(n392), .ZN(n535) );
  INV_X1 U471 ( .A(KEYINPUT1), .ZN(n392) );
  XNOR2_X2 U472 ( .A(n427), .B(G469), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n394), .B(n478), .ZN(n482) );
  XNOR2_X2 U474 ( .A(n464), .B(G116), .ZN(n394) );
  XNOR2_X1 U475 ( .A(n394), .B(n468), .ZN(n474) );
  NAND2_X1 U476 ( .A1(n395), .A2(n348), .ZN(n526) );
  NAND2_X1 U477 ( .A1(n624), .A2(n402), .ZN(n397) );
  XNOR2_X2 U478 ( .A(G119), .B(G113), .ZN(n413) );
  AND2_X1 U479 ( .A1(n450), .A2(n569), .ZN(n403) );
  XOR2_X1 U480 ( .A(KEYINPUT108), .B(n615), .Z(n404) );
  XOR2_X1 U481 ( .A(n420), .B(KEYINPUT30), .Z(n405) );
  NOR2_X1 U482 ( .A1(n710), .A2(n709), .ZN(n406) );
  OR2_X2 U483 ( .A1(n673), .A2(n590), .ZN(n591) );
  XNOR2_X1 U484 ( .A(KEYINPUT69), .B(n574), .ZN(n580) );
  XNOR2_X1 U485 ( .A(n553), .B(n552), .ZN(n559) );
  XNOR2_X1 U486 ( .A(n407), .B(KEYINPUT65), .ZN(n408) );
  XNOR2_X2 U487 ( .A(n472), .B(n408), .ZN(n744) );
  XNOR2_X1 U488 ( .A(KEYINPUT67), .B(G101), .ZN(n409) );
  XNOR2_X1 U489 ( .A(G137), .B(G134), .ZN(n410) );
  XNOR2_X1 U490 ( .A(n410), .B(G131), .ZN(n740) );
  XNOR2_X1 U491 ( .A(n740), .B(G146), .ZN(n411) );
  XNOR2_X2 U492 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n412) );
  NOR2_X1 U493 ( .A1(G953), .A2(G237), .ZN(n456) );
  NAND2_X1 U494 ( .A1(n456), .A2(G210), .ZN(n415) );
  XNOR2_X1 U495 ( .A(G116), .B(KEYINPUT5), .ZN(n414) );
  XNOR2_X1 U496 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U497 ( .A(n478), .B(n416), .ZN(n417) );
  XNOR2_X1 U498 ( .A(n426), .B(n417), .ZN(n641) );
  XNOR2_X1 U499 ( .A(G472), .B(KEYINPUT93), .ZN(n418) );
  XNOR2_X2 U500 ( .A(n536), .B(KEYINPUT103), .ZN(n581) );
  INV_X1 U501 ( .A(G902), .ZN(n475) );
  INV_X1 U502 ( .A(G237), .ZN(n419) );
  NAND2_X1 U503 ( .A1(n475), .A2(n419), .ZN(n491) );
  AND2_X1 U504 ( .A1(n491), .A2(G214), .ZN(n501) );
  INV_X1 U505 ( .A(n501), .ZN(n700) );
  NAND2_X1 U506 ( .A1(n581), .A2(n700), .ZN(n420) );
  XNOR2_X1 U507 ( .A(G107), .B(KEYINPUT89), .ZN(n421) );
  XNOR2_X1 U508 ( .A(n480), .B(n421), .ZN(n424) );
  NAND2_X1 U509 ( .A1(G227), .A2(n731), .ZN(n422) );
  XNOR2_X1 U510 ( .A(n422), .B(G140), .ZN(n423) );
  XNOR2_X1 U511 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U512 ( .A(n426), .B(n425), .ZN(n627) );
  XNOR2_X1 U513 ( .A(n428), .B(KEYINPUT24), .ZN(n429) );
  XOR2_X1 U514 ( .A(KEYINPUT23), .B(n429), .Z(n436) );
  XOR2_X1 U515 ( .A(G110), .B(G137), .Z(n431) );
  NAND2_X1 U516 ( .A1(n731), .A2(G234), .ZN(n433) );
  XNOR2_X1 U517 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n432) );
  XNOR2_X1 U518 ( .A(n433), .B(n432), .ZN(n465) );
  NAND2_X1 U519 ( .A1(G221), .A2(n465), .ZN(n434) );
  INV_X1 U520 ( .A(G125), .ZN(n681) );
  XNOR2_X1 U521 ( .A(n681), .B(G146), .ZN(n486) );
  NAND2_X1 U522 ( .A1(n635), .A2(n475), .ZN(n441) );
  XOR2_X1 U523 ( .A(KEYINPUT74), .B(KEYINPUT25), .Z(n439) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n621) );
  NAND2_X1 U525 ( .A1(n621), .A2(G234), .ZN(n437) );
  XNOR2_X1 U526 ( .A(n437), .B(KEYINPUT20), .ZN(n442) );
  NAND2_X1 U527 ( .A1(n442), .A2(G217), .ZN(n438) );
  XNOR2_X1 U528 ( .A(n439), .B(n438), .ZN(n440) );
  AND2_X1 U529 ( .A1(n442), .A2(G221), .ZN(n444) );
  XNOR2_X1 U530 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n443) );
  XNOR2_X1 U531 ( .A(n444), .B(n443), .ZN(n573) );
  XNOR2_X1 U532 ( .A(n539), .B(KEYINPUT109), .ZN(n450) );
  NAND2_X1 U533 ( .A1(G234), .A2(G237), .ZN(n445) );
  XNOR2_X1 U534 ( .A(n445), .B(KEYINPUT14), .ZN(n448) );
  AND2_X1 U535 ( .A1(G953), .A2(n448), .ZN(n446) );
  NAND2_X1 U536 ( .A1(G902), .A2(n446), .ZN(n505) );
  XNOR2_X1 U537 ( .A(KEYINPUT106), .B(n505), .ZN(n447) );
  NOR2_X1 U538 ( .A1(G900), .A2(n447), .ZN(n449) );
  NAND2_X1 U539 ( .A1(G952), .A2(n448), .ZN(n714) );
  NOR2_X1 U540 ( .A1(G953), .A2(n714), .ZN(n507) );
  OR2_X1 U541 ( .A1(n449), .A2(n507), .ZN(n569) );
  NAND2_X1 U542 ( .A1(n405), .A2(n403), .ZN(n498) );
  XOR2_X1 U543 ( .A(KEYINPUT12), .B(G104), .Z(n452) );
  XNOR2_X1 U544 ( .A(G113), .B(G122), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n452), .B(n451), .ZN(n454) );
  INV_X1 U546 ( .A(KEYINPUT95), .ZN(n453) );
  XNOR2_X1 U547 ( .A(G131), .B(KEYINPUT94), .ZN(n455) );
  XNOR2_X1 U548 ( .A(G143), .B(KEYINPUT97), .ZN(n458) );
  AND2_X1 U549 ( .A1(n456), .A2(G214), .ZN(n457) );
  XNOR2_X1 U550 ( .A(n458), .B(n457), .ZN(n460) );
  XOR2_X1 U551 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n459) );
  XOR2_X1 U552 ( .A(n460), .B(n459), .Z(n461) );
  NAND2_X1 U553 ( .A1(n656), .A2(n475), .ZN(n463) );
  XNOR2_X1 U554 ( .A(KEYINPUT13), .B(G475), .ZN(n462) );
  XNOR2_X2 U555 ( .A(G107), .B(G122), .ZN(n464) );
  NAND2_X1 U556 ( .A1(G217), .A2(n465), .ZN(n467) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n466) );
  XNOR2_X1 U558 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U559 ( .A(KEYINPUT7), .B(KEYINPUT98), .Z(n470) );
  XNOR2_X1 U560 ( .A(G134), .B(KEYINPUT100), .ZN(n469) );
  XNOR2_X1 U561 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U562 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U563 ( .A(n474), .B(n473), .ZN(n724) );
  NAND2_X1 U564 ( .A1(n724), .A2(n475), .ZN(n477) );
  INV_X1 U565 ( .A(G478), .ZN(n476) );
  XNOR2_X1 U566 ( .A(n477), .B(n476), .ZN(n514) );
  XNOR2_X1 U567 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U568 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U569 ( .A(n482), .B(n481), .ZN(n727) );
  NAND2_X1 U570 ( .A1(n731), .A2(G224), .ZN(n483) );
  XNOR2_X1 U571 ( .A(n483), .B(KEYINPUT86), .ZN(n485) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n484) );
  XNOR2_X1 U573 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U574 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U575 ( .A(n727), .B(n488), .ZN(n490) );
  XNOR2_X1 U576 ( .A(n490), .B(n489), .ZN(n648) );
  INV_X1 U577 ( .A(n621), .ZN(n622) );
  OR2_X2 U578 ( .A1(n648), .A2(n622), .ZN(n493) );
  NAND2_X1 U579 ( .A1(n491), .A2(G210), .ZN(n492) );
  XNOR2_X2 U580 ( .A(n493), .B(n492), .ZN(n502) );
  BUF_X1 U581 ( .A(n502), .Z(n494) );
  INV_X1 U582 ( .A(n494), .ZN(n495) );
  NAND2_X1 U583 ( .A1(n346), .A2(n495), .ZN(n496) );
  OR2_X1 U584 ( .A1(n498), .A2(n496), .ZN(n593) );
  XNOR2_X1 U585 ( .A(n593), .B(G143), .ZN(G45) );
  INV_X1 U586 ( .A(KEYINPUT38), .ZN(n497) );
  XNOR2_X1 U587 ( .A(n494), .B(n497), .ZN(n605) );
  OR2_X2 U588 ( .A1(n498), .A2(n605), .ZN(n499) );
  XNOR2_X2 U589 ( .A(n499), .B(KEYINPUT39), .ZN(n602) );
  INV_X1 U590 ( .A(n514), .ZN(n542) );
  AND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n677) );
  NAND2_X1 U592 ( .A1(n602), .A2(n677), .ZN(n618) );
  XOR2_X1 U593 ( .A(G134), .B(KEYINPUT115), .Z(n500) );
  XNOR2_X1 U594 ( .A(n618), .B(n500), .ZN(G36) );
  NOR2_X2 U595 ( .A1(n502), .A2(n501), .ZN(n504) );
  INV_X1 U596 ( .A(KEYINPUT73), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n504), .B(n349), .ZN(n584) );
  NOR2_X1 U598 ( .A1(G898), .A2(n505), .ZN(n506) );
  XOR2_X1 U599 ( .A(KEYINPUT87), .B(n506), .Z(n508) );
  NOR2_X1 U600 ( .A1(n508), .A2(n507), .ZN(n510) );
  INV_X1 U601 ( .A(KEYINPUT88), .ZN(n509) );
  XNOR2_X1 U602 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U603 ( .A1(n584), .A2(n511), .ZN(n513) );
  XNOR2_X1 U604 ( .A(KEYINPUT84), .B(KEYINPUT0), .ZN(n512) );
  INV_X1 U605 ( .A(n534), .ZN(n518) );
  NAND2_X1 U606 ( .A1(n543), .A2(n514), .ZN(n516) );
  INV_X1 U607 ( .A(KEYINPUT101), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n703) );
  INV_X1 U609 ( .A(n573), .ZN(n686) );
  NAND2_X1 U610 ( .A1(n518), .A2(n517), .ZN(n519) );
  INV_X1 U611 ( .A(KEYINPUT102), .ZN(n521) );
  XNOR2_X1 U612 ( .A(n571), .B(n521), .ZN(n687) );
  INV_X1 U613 ( .A(n687), .ZN(n522) );
  AND2_X1 U614 ( .A1(n575), .A2(n522), .ZN(n523) );
  XNOR2_X1 U615 ( .A(G101), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U616 ( .A(n546), .B(n524), .ZN(G3) );
  AND2_X1 U617 ( .A1(n578), .A2(n687), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n526), .B(KEYINPUT32), .ZN(n533) );
  XNOR2_X1 U619 ( .A(n533), .B(G119), .ZN(G21) );
  INV_X1 U620 ( .A(KEYINPUT104), .ZN(n527) );
  XNOR2_X1 U621 ( .A(n528), .B(n527), .ZN(n532) );
  INV_X1 U622 ( .A(n581), .ZN(n530) );
  INV_X1 U623 ( .A(n571), .ZN(n529) );
  AND2_X1 U624 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U625 ( .A1(n532), .A2(n531), .ZN(n663) );
  NAND2_X1 U626 ( .A1(n663), .A2(n533), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n563), .A2(KEYINPUT44), .ZN(n548) );
  BUF_X2 U628 ( .A(n534), .Z(n550) );
  OR2_X1 U629 ( .A1(n536), .A2(n692), .ZN(n537) );
  OR2_X1 U630 ( .A1(n535), .A2(n537), .ZN(n696) );
  OR2_X2 U631 ( .A1(n550), .A2(n696), .ZN(n538) );
  INV_X1 U632 ( .A(n550), .ZN(n541) );
  INV_X1 U633 ( .A(n536), .ZN(n689) );
  NOR2_X1 U634 ( .A1(n539), .A2(n689), .ZN(n540) );
  AND2_X1 U635 ( .A1(n541), .A2(n540), .ZN(n666) );
  INV_X1 U636 ( .A(n677), .ZN(n544) );
  OR2_X1 U637 ( .A1(n543), .A2(n542), .ZN(n600) );
  AND2_X1 U638 ( .A1(n544), .A2(n600), .ZN(n705) );
  INV_X1 U639 ( .A(n705), .ZN(n545) );
  XNOR2_X1 U640 ( .A(KEYINPUT85), .B(KEYINPUT33), .ZN(n549) );
  INV_X1 U641 ( .A(KEYINPUT81), .ZN(n551) );
  XNOR2_X1 U642 ( .A(n551), .B(KEYINPUT35), .ZN(n552) );
  NAND2_X1 U643 ( .A1(n559), .A2(KEYINPUT44), .ZN(n555) );
  INV_X1 U644 ( .A(KEYINPUT83), .ZN(n554) );
  XNOR2_X1 U645 ( .A(n555), .B(n554), .ZN(n556) );
  INV_X1 U646 ( .A(KEYINPUT82), .ZN(n558) );
  BUF_X1 U647 ( .A(n559), .Z(n560) );
  INV_X1 U648 ( .A(n560), .ZN(n562) );
  INV_X1 U649 ( .A(KEYINPUT44), .ZN(n561) );
  AND2_X1 U650 ( .A1(n562), .A2(n561), .ZN(n566) );
  BUF_X1 U651 ( .A(n563), .Z(n564) );
  INV_X1 U652 ( .A(n564), .ZN(n565) );
  NAND2_X1 U653 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U654 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n568) );
  INV_X1 U655 ( .A(n569), .ZN(n570) );
  NOR2_X1 U656 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U657 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U658 ( .A1(n576), .A2(n700), .ZN(n615) );
  NOR2_X1 U659 ( .A1(n615), .A2(n494), .ZN(n577) );
  XNOR2_X1 U660 ( .A(n577), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n579), .A2(n578), .ZN(n680) );
  NAND2_X1 U662 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U663 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n582) );
  BUF_X1 U664 ( .A(n584), .Z(n585) );
  INV_X1 U665 ( .A(n585), .ZN(n586) );
  NOR2_X1 U666 ( .A1(n705), .A2(KEYINPUT47), .ZN(n587) );
  XNOR2_X1 U667 ( .A(n587), .B(KEYINPUT72), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n673), .A2(n588), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n680), .A2(n589), .ZN(n599) );
  INV_X1 U670 ( .A(KEYINPUT47), .ZN(n590) );
  XNOR2_X1 U671 ( .A(n591), .B(KEYINPUT78), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n705), .A2(KEYINPUT47), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U674 ( .A(n594), .B(KEYINPUT75), .ZN(n595) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT77), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n612) );
  INV_X1 U677 ( .A(n600), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n604) );
  INV_X1 U679 ( .A(KEYINPUT40), .ZN(n603) );
  XNOR2_X2 U680 ( .A(n604), .B(n603), .ZN(n662) );
  NAND2_X1 U681 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U682 ( .A1(n704), .A2(n703), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(KEYINPUT41), .ZN(n715) );
  OR2_X1 U684 ( .A1(n715), .A2(n607), .ZN(n609) );
  INV_X1 U685 ( .A(KEYINPUT42), .ZN(n608) );
  NOR2_X2 U686 ( .A1(n662), .A2(n753), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT46), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U689 ( .A(KEYINPUT48), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n614), .B(n613), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n404), .A2(n535), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT43), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n617), .A2(n494), .ZN(n683) );
  AND2_X1 U694 ( .A1(n683), .A2(n618), .ZN(n619) );
  AND2_X1 U695 ( .A1(n622), .A2(KEYINPUT2), .ZN(n623) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n685) );
  NAND2_X1 U697 ( .A1(n722), .A2(G469), .ZN(n629) );
  XNOR2_X1 U698 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n625) );
  XOR2_X1 U699 ( .A(n625), .B(KEYINPUT58), .Z(n626) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n631) );
  INV_X1 U701 ( .A(G952), .ZN(n630) );
  NOR2_X2 U702 ( .A1(n631), .A2(n726), .ZN(n633) );
  INV_X1 U703 ( .A(KEYINPUT121), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(G54) );
  NAND2_X1 U705 ( .A1(n722), .A2(G217), .ZN(n637) );
  XNOR2_X1 U706 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X2 U708 ( .A1(n638), .A2(n726), .ZN(n640) );
  INV_X1 U709 ( .A(KEYINPUT125), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G66) );
  NAND2_X1 U711 ( .A1(n722), .A2(G472), .ZN(n644) );
  BUF_X1 U712 ( .A(n641), .Z(n642) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U714 ( .A1(n645), .A2(n726), .ZN(n647) );
  XNOR2_X1 U715 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G57) );
  NAND2_X1 U717 ( .A1(n722), .A2(G210), .ZN(n653) );
  BUF_X1 U718 ( .A(n648), .Z(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT76), .B(KEYINPUT54), .ZN(n649) );
  XOR2_X1 U720 ( .A(n649), .B(KEYINPUT55), .Z(n650) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X2 U722 ( .A1(n654), .A2(n726), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U724 ( .A1(n722), .A2(G475), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X2 U726 ( .A1(n659), .A2(n726), .ZN(n661) );
  XNOR2_X1 U727 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(G60) );
  XOR2_X1 U729 ( .A(n662), .B(G131), .Z(G33) );
  XNOR2_X1 U730 ( .A(n343), .B(G110), .ZN(G12) );
  XOR2_X1 U731 ( .A(n560), .B(G122), .Z(G24) );
  XOR2_X1 U732 ( .A(G104), .B(KEYINPUT113), .Z(n665) );
  NAND2_X1 U733 ( .A1(n666), .A2(n675), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(G6) );
  XOR2_X1 U735 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n668) );
  NAND2_X1 U736 ( .A1(n666), .A2(n677), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(G107), .B(n669), .ZN(G9) );
  XOR2_X1 U739 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U740 ( .A1(n673), .A2(n677), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(G128), .B(n672), .ZN(G30) );
  NAND2_X1 U743 ( .A1(n673), .A2(n675), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(G146), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n678), .A2(n675), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n676), .B(G113), .ZN(G15) );
  NAND2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n679), .B(G116), .ZN(G18) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U751 ( .A(n683), .B(G140), .ZN(n684) );
  XNOR2_X1 U752 ( .A(KEYINPUT116), .B(n684), .ZN(G42) );
  XNOR2_X1 U753 ( .A(n351), .B(n685), .ZN(n719) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(KEYINPUT49), .B(n688), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U757 ( .A(KEYINPUT117), .B(n691), .Z(n695) );
  NAND2_X1 U758 ( .A1(n535), .A2(n692), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT50), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n697) );
  AND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U762 ( .A(KEYINPUT51), .B(n698), .Z(n699) );
  NOR2_X1 U763 ( .A1(n715), .A2(n699), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n706), .B(KEYINPUT118), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n406), .ZN(n712) );
  XNOR2_X1 U770 ( .A(n712), .B(KEYINPUT52), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n715), .A2(n709), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U774 ( .A1(G953), .A2(n720), .ZN(n721) );
  XNOR2_X1 U775 ( .A(KEYINPUT53), .B(n721), .ZN(G75) );
  NAND2_X1 U776 ( .A1(n722), .A2(G478), .ZN(n723) );
  XOR2_X1 U777 ( .A(n724), .B(n723), .Z(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(G63) );
  BUF_X1 U779 ( .A(n727), .Z(n728) );
  XOR2_X1 U780 ( .A(n728), .B(G101), .Z(n730) );
  NOR2_X1 U781 ( .A1(G898), .A2(n731), .ZN(n729) );
  NOR2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n739) );
  NAND2_X1 U783 ( .A1(n344), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(KEYINPUT126), .ZN(n737) );
  NAND2_X1 U785 ( .A1(G953), .A2(G224), .ZN(n734) );
  XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n734), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(G898), .ZN(n736) );
  NAND2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n739), .B(n738), .ZN(G69) );
  INV_X1 U790 ( .A(n740), .ZN(n741) );
  XNOR2_X1 U791 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n744), .B(n743), .ZN(n748) );
  XNOR2_X1 U793 ( .A(n745), .B(n748), .ZN(n746) );
  NOR2_X1 U794 ( .A1(n746), .A2(G953), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n747), .B(KEYINPUT127), .ZN(n752) );
  XNOR2_X1 U796 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G953), .ZN(n751) );
  NAND2_X1 U799 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U800 ( .A(G137), .B(n753), .Z(G39) );
endmodule

