//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .A3(G137), .ZN(new_n475));
  OAI211_X1 g050(.A(G137), .B(new_n469), .C1(new_n464), .C2(new_n465), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n474), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n474), .A2(new_n496), .A3(G138), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n469), .C1(new_n464), .C2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n501), .A3(KEYINPUT6), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n506), .ZN(new_n514));
  INV_X1    g089(.A(new_n502), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(new_n501), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n513), .A2(new_n519), .A3(new_n521), .ZN(G166));
  XNOR2_X1  g097(.A(KEYINPUT71), .B(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n510), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n512), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n518), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n501), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n501), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n507), .A2(G43), .A3(G543), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n511), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  AND2_X1   g127(.A1(G53), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AND4_X1   g131(.A1(new_n514), .A2(new_n515), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(new_n507), .B2(new_n553), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT74), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n514), .A2(new_n515), .A3(new_n553), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(new_n555), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n507), .A2(new_n553), .A3(new_n556), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g140(.A(KEYINPUT76), .B(G65), .Z(new_n566));
  AND3_X1   g141(.A1(new_n508), .A2(KEYINPUT75), .A3(new_n509), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT75), .B1(new_n508), .B2(new_n509), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G91), .B2(new_n512), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n565), .A2(KEYINPUT77), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT77), .B1(new_n565), .B2(new_n572), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(G299));
  NAND3_X1  g150(.A1(new_n513), .A2(new_n519), .A3(new_n521), .ZN(G303));
  NAND2_X1  g151(.A1(new_n512), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n518), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT78), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n508), .B2(new_n509), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n507), .A2(G86), .A3(new_n510), .ZN(new_n586));
  AND2_X1   g161(.A1(G48), .A2(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n514), .A2(new_n515), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n501), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n507), .A2(G47), .A3(G543), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n511), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  INV_X1    g175(.A(new_n568), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n508), .A2(KEYINPUT75), .A3(new_n509), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G79), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n517), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT80), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(G66), .B1(new_n567), .B2(new_n568), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(new_n604), .C2(new_n517), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n609), .A3(G651), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n514), .A2(G92), .A3(new_n515), .A4(new_n510), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(new_n614), .B1(G54), .B2(new_n518), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n599), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n599), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G280));
  XNOR2_X1  g196(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n546), .A2(new_n619), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n610), .A2(new_n615), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(new_n619), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n472), .A2(new_n473), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n470), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n474), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n487), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n469), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(new_n637), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT83), .Z(G156));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT88), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT87), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT86), .B(G2438), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT85), .ZN(new_n663));
  XOR2_X1   g238(.A(G2451), .B(G2454), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n635), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n673), .B2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n643), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n685), .A3(KEYINPUT89), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n687), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n683), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  NAND2_X1  g277(.A1(G166), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G16), .B2(G22), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(G1971), .C1(G16), .C2(G22), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G23), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G288), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n706), .B(new_n707), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(G6), .ZN(new_n713));
  INV_X1    g288(.A(G305), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT32), .B(G1981), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(new_n711), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n708), .A2(G24), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n708), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n720), .A2(new_n722), .B1(G1986), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n474), .A2(G131), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n487), .A2(G119), .ZN(new_n731));
  OR2_X1    g306(.A1(G95), .A2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n729), .B1(new_n735), .B2(new_n728), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  XOR2_X1   g312(.A(new_n736), .B(new_n737), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n712), .A2(new_n719), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n721), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n726), .A2(G1986), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n727), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(KEYINPUT36), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n727), .A2(new_n744), .A3(new_n740), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n708), .A2(G20), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT23), .Z(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G299), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1956), .ZN(new_n750));
  INV_X1    g325(.A(G19), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n751), .A2(KEYINPUT93), .A3(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT93), .B1(new_n751), .B2(G16), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n547), .C2(new_n708), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n728), .B1(new_n757), .B2(G28), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n756), .B1(new_n758), .B2(new_n759), .C1(new_n642), .C2(new_n728), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n728), .A2(G32), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n487), .A2(G129), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n761), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n760), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n728), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n728), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT29), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n770), .B1(new_n767), .B2(new_n769), .C1(new_n773), .C2(G2090), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G33), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT94), .Z(new_n776));
  AND2_X1   g351(.A1(new_n631), .A2(G127), .ZN(new_n777));
  AND2_X1   g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  OAI21_X1  g353(.A(G2105), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n474), .A2(G139), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT25), .Z(new_n782));
  NAND3_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(new_n728), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2072), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n728), .A2(G26), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT28), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n474), .A2(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n487), .A2(G128), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n728), .A2(G27), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT98), .Z(new_n796));
  AND2_X1   g371(.A1(new_n491), .A2(new_n494), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n496), .B1(new_n474), .B2(G138), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n796), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n785), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n708), .A2(G21), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G286), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G1966), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  NOR4_X1   g383(.A1(new_n755), .A2(new_n774), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G4), .A2(G16), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n616), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT92), .ZN(new_n812));
  INV_X1    g387(.A(G1348), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n708), .A2(G5), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G171), .B2(new_n708), .ZN(new_n816));
  INV_X1    g391(.A(G1961), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G34), .ZN(new_n819));
  AOI21_X1  g394(.A(G29), .B1(new_n819), .B2(KEYINPUT24), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT24), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n480), .B2(new_n728), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2084), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n805), .A2(new_n806), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT96), .Z(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  INV_X1    g402(.A(new_n773), .ZN(new_n828));
  INV_X1    g403(.A(G2090), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n773), .A2(KEYINPUT99), .A3(G2090), .ZN(new_n831));
  AOI211_X1 g406(.A(new_n824), .B(new_n826), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  AND4_X1   g407(.A1(new_n750), .A2(new_n809), .A3(new_n814), .A4(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n746), .A2(new_n833), .ZN(G311));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n746), .A2(new_n835), .A3(new_n833), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n746), .B2(new_n833), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(G150));
  NAND3_X1  g413(.A1(new_n507), .A2(G55), .A3(G543), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n507), .A2(G93), .A3(new_n510), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n508), .B2(new_n509), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  AND2_X1   g420(.A1(G80), .A2(G543), .ZN(new_n846));
  OR3_X1    g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(G651), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n848), .A2(G651), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n841), .B1(new_n853), .B2(new_n847), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n546), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n543), .B(KEYINPUT72), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n540), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n616), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  AOI21_X1  g439(.A(G860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n856), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(G145));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n800), .B(new_n792), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n766), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n783), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n474), .A2(G142), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n487), .A2(G130), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n469), .A2(G118), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n875), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n633), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n735), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n873), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n874), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n873), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n480), .B(new_n642), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n489), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n870), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(new_n887), .B2(new_n884), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT40), .Z(G395));
  XOR2_X1   g465(.A(new_n860), .B(new_n627), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n565), .A2(new_n572), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT77), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n565), .A2(new_n572), .A3(KEYINPUT77), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n616), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n626), .B1(new_n573), .B2(new_n574), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT104), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n891), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT41), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(KEYINPUT105), .B(new_n626), .C1(new_n573), .C2(new_n574), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n896), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n904), .B1(new_n891), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  OAI221_X1 g490(.A(new_n904), .B1(new_n915), .B2(KEYINPUT42), .C1(new_n891), .C2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(G290), .A2(new_n714), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n594), .B(new_n595), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(G305), .A3(new_n591), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G166), .B(G288), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G303), .B(G288), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n919), .A3(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(new_n915), .B2(KEYINPUT42), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n914), .A2(new_n916), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n914), .B2(new_n916), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n856), .A2(new_n619), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  XNOR2_X1  g507(.A(G301), .B(G286), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n852), .A2(new_n855), .B1(new_n858), .B2(new_n540), .ZN(new_n935));
  INV_X1    g510(.A(new_n859), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n857), .A2(new_n859), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n897), .B2(new_n899), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n940), .B(new_n925), .C1(new_n911), .C2(new_n939), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n941), .A2(new_n870), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT107), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n922), .B2(new_n924), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n900), .A2(new_n939), .A3(new_n902), .ZN(new_n948));
  AND4_X1   g523(.A1(KEYINPUT41), .A2(new_n907), .A3(new_n896), .A4(new_n908), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n910), .B1(new_n897), .B2(new_n899), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n938), .A3(new_n937), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n941), .A3(new_n944), .A4(new_n870), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n940), .B1(new_n911), .B2(new_n939), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n947), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n941), .A2(new_n870), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n947), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT43), .B1(new_n942), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n966), .ZN(G397));
  NAND3_X1  g542(.A1(new_n471), .A2(G40), .A3(new_n479), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G164), .B2(G1384), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n800), .A2(KEYINPUT111), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G8), .ZN(new_n975));
  INV_X1    g550(.A(G1976), .ZN(new_n976));
  NOR2_X1   g551(.A1(G288), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT52), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g553(.A1(G288), .A2(new_n976), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT52), .B1(G288), .B2(new_n976), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n974), .A4(G8), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT112), .B(G1981), .Z(new_n983));
  AND4_X1   g558(.A1(new_n586), .A2(new_n585), .A3(new_n588), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT113), .B(G86), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n514), .A2(new_n515), .A3(new_n510), .A4(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n987), .A2(KEYINPUT114), .A3(new_n588), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT114), .B1(new_n987), .B2(new_n588), .ZN(new_n989));
  INV_X1    g564(.A(new_n585), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT49), .B(new_n985), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n987), .A2(new_n588), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n987), .A2(KEYINPUT114), .A3(new_n588), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n585), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G1981), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(KEYINPUT115), .A3(KEYINPUT49), .A4(new_n985), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n995), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT49), .B1(new_n1001), .B2(new_n985), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n975), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(KEYINPUT116), .A3(new_n1005), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n982), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n800), .A2(new_n972), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n968), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n497), .A2(new_n499), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1384), .B1(new_n1014), .B2(new_n797), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(KEYINPUT45), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n800), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT109), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT110), .B(G1971), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n971), .A2(new_n973), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1024), .A2(new_n829), .A3(new_n969), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G166), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1027), .A2(new_n1033), .A3(G8), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1023), .B1(new_n971), .B2(new_n973), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n969), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n829), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1022), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1033), .B1(new_n1041), .B2(G8), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1013), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1044));
  INV_X1    g619(.A(G2078), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1013), .A2(new_n1046), .A3(new_n1019), .A4(new_n1017), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1044), .A2(new_n1045), .B1(new_n1047), .B2(KEYINPUT53), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR4_X1   g624(.A1(new_n1020), .A2(new_n1046), .A3(new_n1049), .A4(G2078), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1024), .A2(new_n969), .A3(new_n1025), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1052), .A2(KEYINPUT124), .A3(new_n817), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT124), .B1(new_n1052), .B2(new_n817), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1049), .B1(new_n1020), .B2(G2078), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1052), .A2(new_n817), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n971), .B2(new_n973), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n969), .A2(new_n1018), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1045), .A2(KEYINPUT53), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1057), .B(new_n1058), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n1063), .B2(G171), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1010), .B(new_n1043), .C1(new_n1056), .C2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1066));
  NAND3_X1  g641(.A1(new_n1051), .A2(G301), .A3(new_n1055), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(G171), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n561), .B2(new_n563), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n572), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1956), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1013), .A2(new_n1017), .A3(new_n1019), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1078), .B2(KEYINPUT121), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1044), .A2(new_n1082), .A3(new_n1077), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1074), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1076), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1052), .A2(new_n813), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n974), .A2(G2067), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n1092), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n616), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1996), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1013), .A2(new_n1098), .A3(new_n1019), .A4(new_n1017), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n974), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n547), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n1092), .A4(new_n626), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1089), .A2(new_n1090), .A3(new_n1097), .A4(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1086), .A2(new_n616), .A3(new_n1093), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1110), .A2(new_n1081), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n968), .A2(G2084), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1024), .A2(new_n1025), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n806), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1024), .A2(new_n1117), .A3(new_n1025), .A4(new_n1113), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(G8), .A3(G286), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1029), .B1(new_n1121), .B2(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G286), .A2(G8), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT122), .Z(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT51), .B(new_n1120), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(G8), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1070), .A2(new_n1112), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n982), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1003), .A2(KEYINPUT116), .A3(new_n1005), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT116), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1029), .B1(new_n1040), .B2(new_n1022), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1034), .B1(new_n1033), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1135), .A2(new_n1137), .A3(new_n1068), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1125), .A2(KEYINPUT62), .A3(new_n1128), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT62), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT126), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1141), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n1139), .A4(new_n1138), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G288), .A2(G1976), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT118), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n984), .B(KEYINPUT117), .Z(new_n1149));
  AOI21_X1  g724(.A(new_n975), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1151));
  NOR2_X1   g726(.A1(new_n1126), .A2(G286), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1041), .A2(G8), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1032), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1035), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1151), .B1(new_n1155), .B2(new_n1135), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1033), .B1(new_n1027), .B2(G8), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1035), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1010), .A3(new_n1152), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1150), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1131), .A2(new_n1142), .A3(new_n1145), .A4(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(G290), .A2(G1986), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n766), .B(new_n1098), .ZN(new_n1164));
  INV_X1    g739(.A(G2067), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n792), .B(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n734), .B(new_n737), .Z(new_n1168));
  NOR2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1163), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n968), .A2(new_n1015), .A3(KEYINPUT45), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1162), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1166), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1175), .B2(new_n766), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1172), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1177), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1172), .B2(new_n1098), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1176), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT47), .Z(new_n1182));
  NOR2_X1   g757(.A1(new_n1169), .A2(new_n1177), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT127), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1163), .A2(new_n1177), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n735), .A2(new_n737), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1167), .A2(new_n1189), .B1(G2067), .B2(new_n792), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1182), .B(new_n1188), .C1(new_n1172), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1174), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g767(.A1(G227), .A2(new_n461), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n668), .A2(new_n701), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1195), .A2(new_n889), .ZN(new_n1196));
  AND2_X1   g770(.A1(new_n1196), .A2(new_n960), .ZN(G308));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n960), .ZN(G225));
endmodule


