//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G116), .ZN(new_n215));
  INV_X1    g0015(.A(G270), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G97), .A2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n217), .B(new_n222), .C1(G58), .C2(G232), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G1), .B2(G20), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n228), .A2(G1), .A3(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G58), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(new_n220), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n213), .B(new_n225), .C1(new_n232), .C2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n216), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n215), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AND3_X1   g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n227), .B2(new_n229), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G50), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n231), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n231), .A2(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(G20), .B2(new_n203), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n258), .B1(G50), .B2(new_n259), .C1(new_n266), .C2(new_n255), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n272), .B1(new_n273), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n263), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n230), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n263), .C2(new_n277), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n256), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n283), .A2(G274), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n284), .A2(new_n281), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n280), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G190), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n280), .A2(new_n286), .A3(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G200), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n267), .A2(new_n268), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n269), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n292), .A2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(new_n290), .A4(new_n269), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n289), .A2(G169), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n267), .B1(new_n291), .B2(G179), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  OAI211_X1 g0106(.A(G226), .B(new_n271), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(G232), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n279), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n287), .A2(G238), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n286), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n315), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n311), .A2(new_n286), .A3(new_n312), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(G179), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n313), .A2(new_n314), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n311), .A2(new_n286), .A3(KEYINPUT13), .A4(new_n312), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G169), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n322), .A2(new_n326), .A3(G169), .A4(new_n323), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n316), .A2(KEYINPUT71), .A3(G179), .A4(new_n318), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n321), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n254), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n230), .A2(G68), .A3(new_n330), .A4(new_n257), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT12), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n259), .B2(G68), .ZN(new_n333));
  INV_X1    g0133(.A(new_n259), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT12), .A3(new_n220), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n331), .A2(new_n338), .A3(new_n333), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n220), .A2(G20), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n341), .B1(new_n261), .B2(new_n273), .C1(new_n202), .C2(new_n264), .ZN(new_n342));
  INV_X1    g0142(.A(new_n255), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT11), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT11), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n329), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n322), .A2(G200), .A3(new_n323), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n316), .A2(G190), .A3(new_n318), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n337), .A2(new_n339), .B1(new_n345), .B2(new_n347), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n357));
  INV_X1    g0157(.A(G107), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n358), .B2(new_n270), .C1(new_n274), .C2(new_n221), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n279), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n287), .A2(G244), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n286), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(G179), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT8), .B(G58), .Z(new_n364));
  NOR2_X1   g0164(.A1(G20), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(KEYINPUT15), .A2(G87), .ZN(new_n367));
  NAND2_X1  g0167(.A1(KEYINPUT15), .A2(G87), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT68), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(KEYINPUT68), .A3(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n366), .B1(new_n231), .B2(new_n273), .C1(new_n373), .C2(new_n261), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n343), .B1(new_n273), .B2(new_n334), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n255), .A2(G77), .A3(new_n257), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G169), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n362), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n363), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n304), .A2(new_n356), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n270), .A2(G257), .A3(new_n271), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n305), .A2(new_n306), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G303), .ZN(new_n385));
  OAI211_X1 g0185(.A(G264), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n279), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT5), .B(G41), .ZN(new_n389));
  INV_X1    g0189(.A(G45), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(G1), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n389), .A2(new_n284), .A3(G274), .A4(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(KEYINPUT5), .A2(G41), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT5), .A2(G41), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(G270), .A3(new_n284), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n259), .A2(G116), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n256), .A2(G33), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n255), .A2(G116), .A3(new_n402), .A4(new_n259), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n263), .A2(G97), .ZN(new_n404));
  AOI21_X1  g0204(.A(G20), .B1(G33), .B2(G283), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n230), .A2(new_n330), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n231), .A2(G116), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT20), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n405), .A2(new_n404), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT20), .ZN(new_n411));
  NOR4_X1   g0211(.A1(new_n255), .A2(new_n410), .A3(new_n411), .A4(new_n407), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n401), .B(new_n403), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n399), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(G169), .A3(new_n397), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT21), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n413), .A2(KEYINPUT21), .A3(G169), .A4(new_n397), .ZN(new_n418));
  INV_X1    g0218(.A(new_n413), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n388), .A2(G190), .A3(new_n392), .A4(new_n396), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n397), .A2(G200), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND4_X1   g0222(.A1(new_n414), .A2(new_n417), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n231), .A2(G107), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT23), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n231), .B(G87), .C1(new_n305), .C2(new_n306), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n427), .A2(KEYINPUT22), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(KEYINPUT22), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n424), .B(new_n426), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n427), .B(KEYINPUT22), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT80), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n424), .A4(new_n426), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(KEYINPUT24), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT24), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(KEYINPUT80), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n343), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(G257), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n439));
  OAI211_X1 g0239(.A(G250), .B(new_n271), .C1(new_n305), .C2(new_n306), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G294), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n279), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n395), .A2(G264), .A3(new_n284), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT83), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n395), .A2(KEYINPUT83), .A3(G264), .A4(new_n284), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n443), .A2(new_n446), .A3(new_n392), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G200), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(new_n444), .A3(new_n392), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(G190), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n334), .B(new_n358), .C1(new_n453), .C2(KEYINPUT25), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT25), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(KEYINPUT81), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n334), .A2(new_n453), .A3(KEYINPUT25), .A4(new_n358), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n255), .A2(new_n402), .A3(new_n259), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n456), .A2(new_n457), .B1(new_n459), .B2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n438), .A2(new_n452), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n438), .A2(new_n460), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n451), .B2(G169), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(G179), .A4(new_n392), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT84), .B1(new_n448), .B2(new_n398), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n451), .A2(new_n463), .A3(G169), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n465), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n423), .A2(new_n461), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n395), .A2(G257), .A3(new_n284), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n392), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n271), .C1(new_n305), .C2(new_n306), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n482), .B2(new_n279), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n449), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n279), .ZN(new_n485));
  INV_X1    g0285(.A(new_n475), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT77), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(KEYINPUT77), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n484), .B1(new_n491), .B2(G190), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT7), .B1(new_n384), .B2(new_n231), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT7), .ZN(new_n494));
  NOR4_X1   g0294(.A1(new_n305), .A2(new_n306), .A3(new_n494), .A4(G20), .ZN(new_n495));
  OAI21_X1  g0295(.A(G107), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT75), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT75), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n498), .B(G107), .C1(new_n493), .C2(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n358), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n358), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n500), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n365), .A2(G77), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n497), .A2(new_n499), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n343), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT76), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n511), .A3(new_n343), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n259), .A2(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n459), .B2(G97), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n492), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n508), .A2(new_n511), .A3(new_n343), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n511), .B1(new_n508), .B2(new_n343), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n488), .B(new_n475), .C1(new_n482), .C2(new_n279), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT77), .B1(new_n485), .B2(new_n486), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n378), .B1(new_n398), .B2(new_n483), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n270), .A2(new_n231), .A3(G68), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n231), .B1(new_n309), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n503), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n309), .B2(G20), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n525), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n343), .B1(new_n373), .B2(new_n334), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n459), .A2(G87), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G238), .B(new_n271), .C1(new_n305), .C2(new_n306), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT78), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT78), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n270), .A2(new_n538), .A3(G238), .A4(new_n271), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G116), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n270), .A2(G244), .A3(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n537), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n279), .ZN(new_n543));
  INV_X1    g0343(.A(new_n391), .ZN(new_n544));
  INV_X1    g0344(.A(G274), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n284), .A2(new_n544), .A3(G250), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n543), .A2(G190), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n535), .B(new_n549), .C1(new_n550), .C2(new_n449), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n459), .A2(KEYINPUT79), .A3(new_n371), .A4(new_n372), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT79), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n458), .B2(new_n373), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n533), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n543), .A2(new_n398), .A3(new_n547), .A4(new_n548), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n550), .C2(G169), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n516), .A2(new_n524), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n260), .B1(new_n255), .B2(new_n257), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n364), .A2(new_n334), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT74), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT73), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G58), .A2(G68), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n231), .B1(new_n234), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n365), .A2(G159), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n566), .ZN(new_n571));
  OAI21_X1  g0371(.A(G20), .B1(new_n571), .B2(new_n201), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(KEYINPUT73), .A3(new_n568), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n495), .ZN(new_n575));
  OR2_X1    g0375(.A1(KEYINPUT3), .A2(G33), .ZN(new_n576));
  NAND2_X1  g0376(.A1(KEYINPUT3), .A2(G33), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(KEYINPUT72), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT72), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n305), .B2(new_n306), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n575), .B1(new_n581), .B2(KEYINPUT7), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n574), .B1(new_n582), .B2(G68), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n255), .B1(new_n583), .B2(KEYINPUT16), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT16), .ZN(new_n585));
  INV_X1    g0385(.A(new_n493), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n220), .B1(new_n586), .B2(new_n575), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n587), .B2(new_n574), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n564), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n270), .A2(G226), .A3(G1698), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n270), .A2(G223), .A3(new_n271), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G87), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n279), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n287), .A2(G232), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n286), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G169), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n594), .A2(G179), .A3(new_n595), .A4(new_n286), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n589), .A2(KEYINPUT18), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT18), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n582), .A2(G68), .ZN(new_n602));
  INV_X1    g0402(.A(new_n574), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(KEYINPUT16), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n343), .A3(new_n588), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n562), .B(KEYINPUT74), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n597), .A2(new_n598), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n596), .A2(new_n449), .ZN(new_n611));
  INV_X1    g0411(.A(G190), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n594), .A2(new_n612), .A3(new_n595), .A4(new_n286), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n614), .A3(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT17), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT17), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n589), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n362), .A2(new_n612), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n362), .A2(G200), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n375), .A4(new_n376), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n610), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NOR4_X1   g0423(.A1(new_n382), .A2(new_n473), .A3(new_n559), .A4(new_n623), .ZN(G372));
  NOR2_X1   g0424(.A1(new_n382), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n551), .A2(new_n557), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT26), .B1(new_n524), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n468), .A2(new_n469), .ZN(new_n628));
  INV_X1    g0428(.A(new_n470), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n464), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n628), .A2(new_n630), .B1(new_n438), .B2(new_n460), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n417), .A2(new_n414), .A3(new_n418), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n461), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n557), .B(new_n627), .C1(new_n559), .C2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n515), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n510), .B2(new_n512), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n491), .A2(G169), .B1(G179), .B2(new_n487), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT85), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n519), .A2(new_n523), .A3(new_n639), .ZN(new_n640));
  AOI211_X1 g0440(.A(KEYINPUT26), .B(new_n626), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n625), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g0443(.A(new_n643), .B(KEYINPUT86), .Z(new_n644));
  AOI22_X1  g0444(.A1(new_n355), .A2(new_n381), .B1(new_n329), .B2(new_n349), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n617), .B1(new_n589), .B2(new_n614), .ZN(new_n646));
  AND4_X1   g0446(.A1(new_n617), .A2(new_n605), .A3(new_n614), .A4(new_n606), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n610), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n302), .B1(new_n649), .B2(new_n299), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT87), .Z(G369));
  NOR2_X1   g0452(.A1(new_n209), .A2(G20), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n256), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n462), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n472), .A2(new_n660), .A3(new_n461), .ZN(new_n661));
  INV_X1    g0461(.A(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n631), .A2(new_n659), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n472), .A2(new_n461), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n419), .A2(new_n662), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n632), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n417), .A2(new_n422), .A3(new_n414), .A4(new_n418), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n666), .A2(new_n663), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n472), .A2(new_n659), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n211), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n529), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n235), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g0484(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n685));
  XNOR2_X1  g0485(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n519), .A2(new_n523), .A3(new_n639), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n639), .B1(new_n519), .B2(new_n523), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n558), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n516), .A2(new_n524), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT89), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n438), .A2(new_n452), .A3(new_n460), .ZN(new_n694));
  INV_X1    g0494(.A(new_n632), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n472), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n692), .A2(new_n693), .A3(new_n558), .A4(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n557), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n524), .A2(new_n626), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT26), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT89), .B1(new_n559), .B2(new_n633), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n691), .A2(new_n697), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n687), .B1(new_n703), .B2(new_n662), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n399), .B1(new_n520), .B2(new_n521), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n550), .A2(new_n466), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n710), .A2(new_n448), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n398), .A3(new_n397), .A4(new_n487), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n491), .A2(KEYINPUT30), .A3(new_n399), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n709), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n659), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n631), .A2(new_n694), .A3(new_n670), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n692), .A2(new_n720), .A3(new_n558), .A4(new_n662), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n705), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n687), .B(new_n662), .C1(new_n634), .C2(new_n641), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n704), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n686), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR2_X1   g0526(.A1(new_n231), .A2(new_n398), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G190), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(KEYINPUT92), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT33), .B(G317), .Z(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(G190), .A3(new_n449), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n231), .A2(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(new_n612), .A3(G200), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(G303), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n738), .A2(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n270), .B1(new_n746), .B2(G329), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n727), .A2(new_n744), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n728), .A2(new_n612), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n743), .B(new_n750), .C1(G326), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n612), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n231), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n737), .B(new_n752), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n751), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n202), .ZN(new_n758));
  INV_X1    g0558(.A(new_n732), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n384), .B1(new_n759), .B2(G68), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n741), .A2(new_n528), .ZN(new_n761));
  INV_X1    g0561(.A(G159), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n745), .A2(KEYINPUT32), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n735), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n761), .B(new_n763), .C1(G58), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n740), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G107), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT32), .B1(new_n745), .B2(new_n762), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n273), .C2(new_n749), .ZN(new_n769));
  INV_X1    g0569(.A(new_n755), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(G97), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n760), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n756), .B1(new_n758), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n230), .B1(G20), .B2(new_n378), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT90), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n249), .A2(G45), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n578), .A2(new_n580), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n679), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n785), .B(new_n788), .C1(G45), .C2(new_n235), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n211), .A2(G355), .A3(new_n270), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(G116), .C2(new_n211), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n773), .A2(new_n778), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n256), .B1(new_n653), .B2(G45), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n680), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n792), .B(new_n795), .C1(new_n671), .C2(new_n782), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT94), .Z(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(new_n671), .B2(G330), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G330), .B2(new_n671), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(G396));
  NAND2_X1  g0600(.A1(new_n642), .A2(new_n662), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n377), .A2(new_n659), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n622), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n380), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n380), .A2(new_n659), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n805), .B1(new_n380), .B2(new_n803), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n662), .B(new_n809), .C1(new_n634), .C2(new_n641), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(new_n722), .ZN(new_n812));
  INV_X1    g0612(.A(new_n795), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n755), .A2(new_n501), .B1(new_n740), .B2(new_n528), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n384), .B1(new_n749), .B2(new_n215), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n759), .C2(G283), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n757), .A2(new_n742), .B1(new_n753), .B2(new_n735), .ZN(new_n818));
  INV_X1    g0618(.A(new_n741), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G107), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(new_n748), .C2(new_n745), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT95), .Z(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n787), .B1(new_n823), .B2(new_n745), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n202), .A2(new_n741), .B1(new_n740), .B2(new_n220), .ZN(new_n825));
  INV_X1    g0625(.A(new_n749), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n764), .A2(G143), .B1(new_n826), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n757), .C1(new_n732), .C2(new_n262), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n824), .B(new_n825), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .C1(new_n233), .C2(new_n755), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n813), .B1(new_n833), .B2(new_n778), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n778), .A2(new_n779), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(G77), .B2(new_n836), .C1(new_n780), .C2(new_n809), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n814), .A2(new_n837), .ZN(G384));
  XOR2_X1   g0638(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n839));
  INV_X1    g0639(.A(new_n657), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n584), .B1(KEYINPUT16), .B2(new_n583), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n560), .B2(new_n561), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT18), .B1(new_n589), .B2(new_n599), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n607), .A2(new_n601), .A3(new_n608), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n840), .B(new_n842), .C1(new_n648), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n597), .A2(new_n598), .A3(new_n657), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n607), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n615), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n842), .A2(new_n847), .B1(new_n589), .B2(new_n614), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n849), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n846), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n846), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n719), .A2(new_n721), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT96), .B1(new_n353), .B2(new_n662), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT96), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n349), .A2(new_n858), .A3(new_n659), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n354), .B(new_n860), .C1(new_n329), .C2(new_n349), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n356), .A2(new_n860), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n807), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n839), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n846), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(new_n847), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n615), .B1(new_n589), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT97), .B1(new_n607), .B2(new_n847), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(new_n849), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n848), .A2(KEYINPUT97), .A3(KEYINPUT37), .A4(new_n615), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n657), .B1(new_n610), .B2(new_n619), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n607), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n867), .B1(new_n875), .B2(KEYINPUT38), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n350), .A2(new_n355), .B1(new_n857), .B2(new_n859), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n809), .B1(new_n877), .B2(new_n861), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n721), .B2(new_n719), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(KEYINPUT40), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n866), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n625), .A2(new_n856), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n881), .B(new_n882), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(G330), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n625), .B1(new_n704), .B2(new_n724), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n650), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n884), .B(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(KEYINPUT98), .B(KEYINPUT100), .Z(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT39), .B1(new_n853), .B2(new_n854), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n867), .C1(new_n875), .C2(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n329), .A2(new_n349), .A3(new_n662), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n877), .A2(new_n861), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n810), .B2(new_n806), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n853), .B2(new_n854), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n845), .A2(new_n657), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n889), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n256), .B2(new_n653), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n215), .B1(new_n505), .B2(KEYINPUT35), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n232), .C1(KEYINPUT35), .C2(new_n505), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n566), .A2(G77), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n235), .A2(new_n908), .B1(G50), .B2(new_n220), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(G1), .A3(new_n209), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n907), .A3(new_n910), .ZN(G367));
  OAI211_X1 g0711(.A(new_n516), .B(new_n524), .C1(new_n636), .C2(new_n662), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n519), .A2(new_n523), .A3(new_n659), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n677), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(KEYINPUT44), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT44), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n677), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n677), .A2(new_n914), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT45), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT45), .B1(new_n677), .B2(new_n914), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n916), .A2(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n667), .B(new_n672), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n725), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n680), .B(KEYINPUT41), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n794), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n914), .A2(KEYINPUT101), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT101), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n912), .A2(new_n913), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n631), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n659), .B1(new_n932), .B2(new_n524), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT43), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n914), .A2(new_n675), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT42), .Z(new_n937));
  NOR2_X1   g0737(.A1(new_n535), .A2(new_n662), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n626), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n698), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n934), .A2(new_n935), .A3(new_n937), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n935), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n936), .B(KEYINPUT42), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n944), .B(new_n945), .C1(new_n933), .C2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n929), .ZN(new_n948));
  INV_X1    g0748(.A(new_n931), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n674), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT103), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT103), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n943), .A2(new_n947), .A3(new_n953), .A4(new_n950), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n950), .B1(new_n943), .B2(new_n947), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT102), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n952), .B(new_n954), .C1(KEYINPUT102), .C2(new_n956), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n928), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(G317), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n786), .B1(new_n961), .B2(new_n745), .C1(new_n732), .C2(new_n753), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G107), .A2(new_n770), .B1(new_n764), .B2(G303), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n766), .A2(G97), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n748), .C2(new_n757), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n741), .A2(new_n215), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n962), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n738), .B2(new_n749), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n749), .A2(new_n202), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n740), .A2(new_n273), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n755), .A2(new_n220), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G150), .C2(new_n764), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n741), .A2(new_n233), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n270), .B1(new_n745), .B2(new_n828), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(G143), .C2(new_n751), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n973), .B(new_n976), .C1(new_n762), .C2(new_n732), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n969), .B1(new_n970), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n813), .B1(new_n979), .B2(new_n778), .ZN(new_n980));
  INV_X1    g0780(.A(new_n788), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n784), .B1(new_n211), .B2(new_n373), .C1(new_n245), .C2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT104), .Z(new_n983));
  OAI211_X1 g0783(.A(new_n980), .B(new_n983), .C1(new_n782), .C2(new_n941), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n960), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(G387));
  OAI22_X1  g0787(.A1(new_n735), .A2(new_n961), .B1(new_n749), .B2(new_n742), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n759), .A2(G311), .B1(KEYINPUT106), .B2(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(KEYINPUT106), .B2(new_n988), .C1(new_n734), .C2(new_n757), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT48), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n738), .B2(new_n755), .C1(new_n753), .C2(new_n741), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT49), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n746), .A2(G326), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n787), .B1(G116), .B2(new_n766), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n786), .B1(G150), .B2(new_n746), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n964), .C1(new_n273), .C2(new_n741), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT105), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n373), .A2(new_n755), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n757), .A2(new_n762), .B1(new_n202), .B2(new_n735), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n759), .C2(new_n364), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1001), .B(new_n1004), .C1(new_n220), .C2(new_n749), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(G116), .B(new_n529), .C1(G68), .C2(G77), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n260), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT50), .B1(new_n260), .B2(G50), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1007), .A2(new_n390), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n981), .B1(new_n241), .B2(G45), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n679), .A2(new_n384), .A3(new_n682), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(G107), .B2(new_n211), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1006), .A2(new_n778), .B1(new_n784), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n661), .A2(new_n664), .A3(new_n783), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n795), .A3(new_n1016), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n704), .A2(new_n925), .A3(new_n724), .A4(new_n722), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n925), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n680), .B1(new_n725), .B2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1017), .B1(new_n793), .B2(new_n925), .C1(new_n1018), .C2(new_n1020), .ZN(G393));
  NAND2_X1  g0821(.A1(new_n923), .A2(new_n673), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n674), .B1(new_n921), .B2(new_n922), .C1(new_n916), .C2(new_n918), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n725), .A2(new_n1019), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(KEYINPUT108), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT108), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1018), .B2(new_n923), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1022), .A2(new_n1023), .B1(new_n725), .B2(new_n1019), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1026), .B(new_n680), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1022), .A2(new_n1023), .A3(new_n794), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n783), .B1(new_n949), .B2(new_n948), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n784), .B1(new_n501), .B2(new_n211), .C1(new_n252), .C2(new_n981), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n787), .B1(new_n260), .B2(new_n749), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n759), .B2(G50), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n757), .A2(new_n262), .B1(new_n762), .B2(new_n735), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n746), .A2(G143), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n740), .A2(new_n528), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n755), .A2(new_n273), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G68), .C2(new_n819), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n270), .B1(new_n746), .B2(G322), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n767), .C1(new_n738), .C2(new_n741), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT107), .Z(new_n1045));
  OAI22_X1  g0845(.A1(new_n757), .A2(new_n961), .B1(new_n748), .B2(new_n735), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n759), .A2(G303), .B1(G294), .B2(new_n826), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n755), .A2(new_n215), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1042), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n813), .B1(new_n1051), .B2(new_n778), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1032), .A2(new_n1033), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1030), .A2(new_n1031), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT109), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1030), .A2(KEYINPUT109), .A3(new_n1031), .A4(new_n1053), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(G390));
  INV_X1    g0858(.A(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n716), .A2(new_n659), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT31), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n559), .A2(new_n473), .A3(new_n659), .ZN(new_n1065));
  OAI211_X1 g0865(.A(G330), .B(new_n809), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n897), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n856), .A2(G330), .A3(new_n864), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1067), .A2(new_n1068), .B1(new_n806), .B2(new_n810), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n703), .A2(new_n662), .A3(new_n804), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1067), .A2(new_n1070), .A3(new_n806), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(KEYINPUT111), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT111), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n879), .A2(new_n1073), .A3(G330), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1069), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n625), .A2(G330), .A3(new_n856), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n885), .A2(new_n650), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1059), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n885), .A2(new_n650), .A3(new_n1077), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n810), .A2(new_n806), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1073), .B1(new_n879), .B2(G330), .ZN(new_n1084));
  AND4_X1   g0884(.A1(new_n1073), .A2(new_n856), .A3(G330), .A4(new_n864), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1067), .A2(new_n1070), .A3(new_n806), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1080), .A2(new_n1088), .A3(KEYINPUT112), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1079), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n897), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1082), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n893), .B1(new_n894), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n894), .B(KEYINPUT110), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n876), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1070), .A2(new_n806), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n1091), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1068), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n890), .B(new_n892), .C1(new_n898), .C2(new_n895), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n897), .B1(new_n1070), .B2(new_n806), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1086), .C1(new_n1100), .C2(new_n1095), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1090), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT113), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1090), .A2(new_n1102), .A3(KEYINPUT113), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1105), .A2(new_n680), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n890), .A2(new_n892), .A3(new_n779), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n759), .A2(G107), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n384), .B1(new_n749), .B2(new_n501), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n761), .B(new_n1113), .C1(G68), .C2(new_n766), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n746), .A2(G294), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n735), .A2(new_n215), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1116), .B(new_n1040), .C1(G283), .C2(new_n751), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n759), .A2(G137), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n741), .A2(new_n262), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n735), .A2(new_n823), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n755), .A2(new_n762), .B1(new_n740), .B2(new_n202), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G128), .C2(new_n751), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n384), .B1(new_n746), .B2(G125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1119), .A2(new_n1122), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n749), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1118), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n778), .B1(new_n260), .B2(new_n835), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1111), .A2(new_n795), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1102), .B2(new_n793), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1110), .A2(new_n1135), .ZN(G378));
  NAND3_X1  g0936(.A1(new_n866), .A2(G330), .A3(new_n880), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n267), .A2(new_n840), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n299), .B2(new_n303), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1138), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1141), .B(new_n302), .C1(new_n295), .C2(new_n298), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT55), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT55), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1145), .A2(KEYINPUT56), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT56), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1137), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n866), .A3(G330), .A4(new_n880), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n902), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n901), .A3(new_n1152), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT117), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT117), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n1157), .A3(new_n902), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n794), .A3(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n759), .A2(G132), .B1(G128), .B2(new_n764), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G150), .A2(new_n770), .B1(new_n751), .B2(G125), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n741), .C2(new_n1129), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G137), .B2(new_n826), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n766), .B2(G159), .ZN(new_n1165));
  XOR2_X1   g0965(.A(KEYINPUT115), .B(G124), .Z(new_n1166));
  AOI21_X1  g0966(.A(G33), .B1(new_n746), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n732), .A2(new_n501), .B1(new_n373), .B2(new_n749), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n972), .B1(G77), .B2(new_n819), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n277), .C1(new_n738), .C2(new_n745), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1169), .A2(new_n787), .A3(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G107), .A2(new_n764), .B1(new_n766), .B2(G58), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n215), .C2(new_n757), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT58), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G41), .B1(new_n787), .B2(G33), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1168), .B(new_n1175), .C1(G50), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n813), .B1(new_n1177), .B2(new_n778), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(G50), .B2(new_n836), .C1(new_n1149), .C2(new_n780), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT116), .Z(new_n1180));
  AND2_X1   g0980(.A1(new_n1159), .A2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1108), .A2(new_n1080), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1080), .A2(new_n1088), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1078), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1154), .A2(KEYINPUT118), .A3(new_n1155), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1153), .A2(new_n902), .A3(KEYINPUT118), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n680), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1181), .B1(new_n1184), .B2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1090), .A2(new_n927), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1091), .A2(new_n780), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n813), .B1(new_n835), .B2(new_n220), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT119), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n732), .A2(new_n215), .B1(new_n358), .B2(new_n749), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT120), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G294), .A2(new_n751), .B1(new_n764), .B2(G283), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n501), .B2(new_n741), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1199), .A2(new_n1002), .A3(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n270), .B(new_n971), .C1(G303), .C2(new_n746), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n746), .A2(G128), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n735), .A2(new_n828), .B1(new_n741), .B2(new_n762), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n751), .A2(G132), .B1(new_n766), .B2(G58), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n786), .B1(G150), .B2(new_n826), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n732), .C2(new_n1129), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1205), .B(new_n1208), .C1(G50), .C2(new_n770), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1202), .A2(new_n1203), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n778), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1197), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT121), .Z(new_n1213));
  OAI22_X1  g1013(.A1(new_n1076), .A2(new_n793), .B1(new_n1195), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1194), .A2(new_n1215), .ZN(G381));
  NOR2_X1   g1016(.A1(G375), .A2(G378), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1217), .A2(new_n986), .A3(new_n1218), .A4(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n658), .A2(G213), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT122), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT123), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(G407), .A2(G213), .A3(new_n1224), .ZN(G409));
  NAND3_X1  g1025(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1078), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1226), .A2(new_n1185), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n681), .B1(new_n1193), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1214), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT124), .B1(new_n1230), .B2(G384), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1080), .A2(new_n1088), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n680), .B1(new_n1232), .B2(KEYINPUT60), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1226), .A2(new_n1185), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1215), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(G384), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1230), .A2(G384), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1231), .A2(new_n1238), .A3(KEYINPUT63), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1078), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1189), .A4(new_n1188), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n680), .A3(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(G378), .A2(new_n1246), .A3(new_n1181), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1183), .A2(new_n927), .A3(new_n1158), .A4(new_n1156), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1188), .A2(new_n1189), .A3(new_n794), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1180), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1135), .A3(new_n1110), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1223), .B(new_n1240), .C1(new_n1247), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n986), .A2(G390), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1056), .B(new_n1057), .C1(new_n960), .C2(new_n985), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  XOR2_X1   g1055(.A(G393), .B(G396), .Z(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(new_n1256), .A3(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1252), .A2(KEYINPUT61), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1231), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1263));
  INV_X1    g1063(.A(G2897), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1222), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1223), .A2(G2897), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1263), .A2(KEYINPUT125), .A3(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1266), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1090), .A2(KEYINPUT113), .A3(new_n1102), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT113), .B1(new_n1090), .B2(new_n1102), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1186), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1134), .B1(new_n1275), .B2(new_n680), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1251), .B1(G375), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1222), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1262), .B1(new_n1272), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1263), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1277), .A2(new_n1222), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1261), .B1(new_n1279), .B2(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1253), .A2(new_n1256), .A3(new_n1254), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1256), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT126), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1258), .A2(new_n1287), .A3(new_n1259), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1223), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1263), .A2(new_n1290), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1281), .A2(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1263), .A2(KEYINPUT125), .A3(new_n1267), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT125), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1294), .B1(new_n1298), .B2(new_n1291), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1289), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1283), .A2(new_n1300), .ZN(G405));
  NAND3_X1  g1101(.A1(G375), .A2(new_n1276), .A3(new_n1263), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1263), .B1(G375), .B2(new_n1276), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1259), .B(new_n1258), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1260), .A2(new_n1306), .A3(new_n1302), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1247), .A2(KEYINPUT127), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


