

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U554 ( .A1(n686), .A2(n798), .ZN(n732) );
  XOR2_X1 U555 ( .A(n732), .B(n687), .Z(n717) );
  NOR2_X1 U556 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  XOR2_X1 U558 ( .A(KEYINPUT32), .B(n744), .Z(n520) );
  INV_X1 U559 ( .A(KEYINPUT64), .ZN(n704) );
  AND2_X1 U560 ( .A1(n688), .A2(n717), .ZN(n690) );
  NOR2_X1 U561 ( .A1(G171), .A2(n699), .ZN(n692) );
  INV_X1 U562 ( .A(n1011), .ZN(n754) );
  NAND2_X1 U563 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U564 ( .A1(n520), .A2(n752), .ZN(n769) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n798) );
  INV_X1 U566 ( .A(KEYINPUT89), .ZN(n532) );
  XNOR2_X1 U567 ( .A(n533), .B(n532), .ZN(n535) );
  AND2_X2 U568 ( .A1(n531), .A2(G2105), .ZN(n889) );
  NOR2_X1 U569 ( .A1(G651), .A2(n647), .ZN(n648) );
  XNOR2_X1 U570 ( .A(KEYINPUT76), .B(n594), .ZN(n1019) );
  NOR2_X1 U571 ( .A1(n543), .A2(n542), .ZN(G164) );
  INV_X1 U572 ( .A(G651), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G543), .A2(n524), .ZN(n521) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n521), .Z(n652) );
  NAND2_X1 U575 ( .A1(G64), .A2(n652), .ZN(n523) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n647) );
  NAND2_X1 U577 ( .A1(G52), .A2(n648), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U580 ( .A1(G90), .A2(n638), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n647), .A2(n524), .ZN(n639) );
  NAND2_X1 U582 ( .A1(G77), .A2(n639), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U584 ( .A(KEYINPUT9), .B(n527), .Z(n528) );
  XNOR2_X1 U585 ( .A(KEYINPUT70), .B(n528), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n530), .A2(n529), .ZN(G171) );
  INV_X1 U587 ( .A(G2104), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n889), .A2(G126), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n890), .A2(G114), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U591 ( .A(KEYINPUT90), .B(n536), .ZN(n543) );
  INV_X1 U592 ( .A(G2105), .ZN(n563) );
  AND2_X1 U593 ( .A1(n563), .A2(G2104), .ZN(n884) );
  NAND2_X1 U594 ( .A1(n884), .A2(G102), .ZN(n541) );
  XNOR2_X1 U595 ( .A(KEYINPUT68), .B(KEYINPUT17), .ZN(n538) );
  NOR2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XNOR2_X1 U597 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U598 ( .A(KEYINPUT67), .B(n539), .ZN(n559) );
  NAND2_X1 U599 ( .A1(G138), .A2(n559), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G85), .A2(n638), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G72), .A2(n639), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G60), .A2(n652), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G47), .A2(n648), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U607 ( .A1(n549), .A2(n548), .ZN(G290) );
  NAND2_X1 U608 ( .A1(G111), .A2(n890), .ZN(n551) );
  BUF_X1 U609 ( .A(n559), .Z(n885) );
  NAND2_X1 U610 ( .A1(G135), .A2(n885), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n889), .A2(G123), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT18), .B(n552), .Z(n553) );
  NOR2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n884), .A2(G99), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n953) );
  XNOR2_X1 U617 ( .A(G2096), .B(n953), .ZN(n557) );
  OR2_X1 U618 ( .A1(G2100), .A2(n557), .ZN(G156) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  INV_X1 U623 ( .A(G57), .ZN(G237) );
  NAND2_X1 U624 ( .A1(G113), .A2(n890), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT66), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n559), .A2(G137), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT69), .B(n560), .Z(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n796) );
  AND2_X1 U629 ( .A1(n563), .A2(G101), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G2104), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT23), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT65), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G125), .A2(n889), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n685) );
  NOR2_X1 U635 ( .A1(n796), .A2(n685), .ZN(G160) );
  NAND2_X1 U636 ( .A1(n639), .A2(G76), .ZN(n569) );
  XNOR2_X1 U637 ( .A(KEYINPUT78), .B(n569), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n638), .A2(G89), .ZN(n570) );
  XNOR2_X1 U639 ( .A(KEYINPUT4), .B(n570), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT5), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G63), .A2(n652), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G51), .A2(n648), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT6), .B(n576), .Z(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U648 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U649 ( .A1(G94), .A2(G452), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U652 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U653 ( .A(G223), .B(KEYINPUT73), .ZN(n832) );
  NAND2_X1 U654 ( .A1(n832), .A2(G567), .ZN(n582) );
  XOR2_X1 U655 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  INV_X1 U656 ( .A(G860), .ZN(n614) );
  NAND2_X1 U657 ( .A1(n638), .A2(G81), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G68), .A2(n639), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(n586), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n588) );
  NAND2_X1 U663 ( .A1(G56), .A2(n652), .ZN(n587) );
  XNOR2_X1 U664 ( .A(n588), .B(n587), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G43), .A2(n648), .ZN(n589) );
  XNOR2_X1 U666 ( .A(KEYINPUT75), .B(n589), .ZN(n590) );
  NOR2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  OR2_X1 U669 ( .A1(n614), .A2(n1019), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G54), .A2(n648), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G92), .A2(n638), .ZN(n596) );
  NAND2_X1 U674 ( .A1(G79), .A2(n639), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G66), .A2(n652), .ZN(n597) );
  XNOR2_X1 U677 ( .A(KEYINPUT77), .B(n597), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n602), .B(KEYINPUT15), .ZN(n903) );
  INV_X1 U681 ( .A(n903), .ZN(n1000) );
  INV_X1 U682 ( .A(G868), .ZN(n665) );
  NAND2_X1 U683 ( .A1(n1000), .A2(n665), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G78), .A2(n639), .ZN(n606) );
  NAND2_X1 U686 ( .A1(G65), .A2(n652), .ZN(n605) );
  NAND2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n638), .A2(G91), .ZN(n607) );
  XOR2_X1 U689 ( .A(KEYINPUT72), .B(n607), .Z(n608) );
  NOR2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n648), .A2(G53), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(G299) );
  NOR2_X1 U693 ( .A1(G286), .A2(n665), .ZN(n613) );
  NOR2_X1 U694 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U695 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U696 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n615), .A2(n903), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U699 ( .A1(n1019), .A2(G868), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G868), .A2(n903), .ZN(n617) );
  NOR2_X1 U701 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U703 ( .A1(G559), .A2(n903), .ZN(n620) );
  XNOR2_X1 U704 ( .A(n620), .B(n1019), .ZN(n662) );
  NOR2_X1 U705 ( .A1(n662), .A2(G860), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G93), .A2(n638), .ZN(n622) );
  NAND2_X1 U707 ( .A1(G67), .A2(n652), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G80), .A2(n639), .ZN(n623) );
  XNOR2_X1 U710 ( .A(KEYINPUT79), .B(n623), .ZN(n624) );
  NOR2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n648), .A2(G55), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n664) );
  XOR2_X1 U714 ( .A(n664), .B(KEYINPUT80), .Z(n628) );
  XNOR2_X1 U715 ( .A(n629), .B(n628), .ZN(G145) );
  NAND2_X1 U716 ( .A1(G86), .A2(n638), .ZN(n631) );
  NAND2_X1 U717 ( .A1(G61), .A2(n652), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n639), .A2(G73), .ZN(n632) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n648), .A2(G48), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G50), .A2(n648), .ZN(n637) );
  XOR2_X1 U725 ( .A(KEYINPUT82), .B(n637), .Z(n644) );
  NAND2_X1 U726 ( .A1(G88), .A2(n638), .ZN(n641) );
  NAND2_X1 U727 ( .A1(G75), .A2(n639), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U729 ( .A(KEYINPUT83), .B(n642), .Z(n643) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n652), .A2(G62), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(G303) );
  INV_X1 U733 ( .A(G303), .ZN(G166) );
  NAND2_X1 U734 ( .A1(n647), .A2(G87), .ZN(n654) );
  NAND2_X1 U735 ( .A1(G49), .A2(n648), .ZN(n650) );
  NAND2_X1 U736 ( .A1(G74), .A2(G651), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U740 ( .A(KEYINPUT81), .B(n655), .Z(G288) );
  INV_X1 U741 ( .A(G299), .ZN(n1009) );
  XNOR2_X1 U742 ( .A(n1009), .B(G305), .ZN(n661) );
  XNOR2_X1 U743 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U744 ( .A(G290), .B(G166), .ZN(n656) );
  XNOR2_X1 U745 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U746 ( .A(n658), .B(G288), .Z(n659) );
  XNOR2_X1 U747 ( .A(n664), .B(n659), .ZN(n660) );
  XNOR2_X1 U748 ( .A(n661), .B(n660), .ZN(n902) );
  XNOR2_X1 U749 ( .A(n662), .B(n902), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U752 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(KEYINPUT20), .ZN(n669) );
  XNOR2_X1 U755 ( .A(n669), .B(KEYINPUT85), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n670), .A2(G2090), .ZN(n671) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(KEYINPUT86), .B(G44), .ZN(n673) );
  XNOR2_X1 U760 ( .A(n673), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G235), .A2(G236), .ZN(n674) );
  XNOR2_X1 U762 ( .A(n674), .B(KEYINPUT87), .ZN(n675) );
  NOR2_X1 U763 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U764 ( .A1(G108), .A2(n676), .ZN(n836) );
  NAND2_X1 U765 ( .A1(n836), .A2(G567), .ZN(n681) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U768 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G96), .A2(n679), .ZN(n837) );
  NAND2_X1 U770 ( .A1(n837), .A2(G2106), .ZN(n680) );
  NAND2_X1 U771 ( .A1(n681), .A2(n680), .ZN(n838) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U773 ( .A1(n838), .A2(n682), .ZN(n835) );
  NAND2_X1 U774 ( .A1(n835), .A2(G36), .ZN(n683) );
  XNOR2_X1 U775 ( .A(KEYINPUT88), .B(n683), .ZN(G176) );
  XNOR2_X1 U776 ( .A(G1981), .B(G305), .ZN(n1006) );
  XOR2_X1 U777 ( .A(G2078), .B(KEYINPUT25), .Z(n926) );
  INV_X1 U778 ( .A(n926), .ZN(n688) );
  INV_X1 U779 ( .A(G40), .ZN(n684) );
  OR2_X1 U780 ( .A1(n685), .A2(n684), .ZN(n795) );
  NOR2_X1 U781 ( .A1(n796), .A2(n795), .ZN(n686) );
  INV_X1 U782 ( .A(KEYINPUT95), .ZN(n687) );
  INV_X1 U783 ( .A(n732), .ZN(n707) );
  NOR2_X1 U784 ( .A1(n707), .A2(G1961), .ZN(n689) );
  NOR2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U786 ( .A(KEYINPUT96), .B(n691), .Z(n699) );
  XNOR2_X1 U787 ( .A(n692), .B(KEYINPUT100), .ZN(n697) );
  NAND2_X1 U788 ( .A1(G8), .A2(n732), .ZN(n774) );
  NOR2_X1 U789 ( .A1(G1966), .A2(n774), .ZN(n751) );
  NOR2_X1 U790 ( .A1(G2084), .A2(n732), .ZN(n747) );
  NOR2_X1 U791 ( .A1(n751), .A2(n747), .ZN(n693) );
  NAND2_X1 U792 ( .A1(G8), .A2(n693), .ZN(n694) );
  XNOR2_X1 U793 ( .A(KEYINPUT30), .B(n694), .ZN(n695) );
  NOR2_X1 U794 ( .A1(n695), .A2(G168), .ZN(n696) );
  NOR2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U796 ( .A(n698), .B(KEYINPUT31), .Z(n745) );
  NAND2_X1 U797 ( .A1(n699), .A2(G171), .ZN(n730) );
  AND2_X1 U798 ( .A1(n707), .A2(G1996), .ZN(n700) );
  XOR2_X1 U799 ( .A(n700), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U800 ( .A1(n732), .A2(G1341), .ZN(n701) );
  NAND2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n1019), .A2(n703), .ZN(n705) );
  XNOR2_X1 U803 ( .A(n705), .B(n704), .ZN(n711) );
  INV_X1 U804 ( .A(G2067), .ZN(n925) );
  INV_X1 U805 ( .A(n717), .ZN(n706) );
  NOR2_X1 U806 ( .A1(n925), .A2(n706), .ZN(n709) );
  INV_X1 U807 ( .A(G1348), .ZN(n999) );
  NOR2_X1 U808 ( .A1(n707), .A2(n999), .ZN(n708) );
  NOR2_X1 U809 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n903), .A2(n712), .ZN(n710) );
  NAND2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n714) );
  OR2_X1 U812 ( .A1(n903), .A2(n712), .ZN(n713) );
  NAND2_X1 U813 ( .A1(n714), .A2(n713), .ZN(n721) );
  XOR2_X1 U814 ( .A(KEYINPUT27), .B(KEYINPUT97), .Z(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(G2072), .ZN(n715) );
  XNOR2_X1 U816 ( .A(n716), .B(n715), .ZN(n719) );
  INV_X1 U817 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U818 ( .A1(n717), .A2(n1008), .ZN(n718) );
  NOR2_X1 U819 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U820 ( .A1(n722), .A2(n1009), .ZN(n720) );
  NAND2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n726) );
  NOR2_X1 U822 ( .A1(n722), .A2(n1009), .ZN(n724) );
  XOR2_X1 U823 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n723) );
  XNOR2_X1 U824 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U825 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U826 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n727) );
  XNOR2_X1 U827 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U828 ( .A1(n730), .A2(n729), .ZN(n746) );
  INV_X1 U829 ( .A(G8), .ZN(n738) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n774), .ZN(n731) );
  XOR2_X1 U831 ( .A(KEYINPUT101), .B(n731), .Z(n734) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U833 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U834 ( .A(n735), .B(KEYINPUT102), .ZN(n736) );
  NAND2_X1 U835 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n740) );
  AND2_X1 U837 ( .A1(n746), .A2(n740), .ZN(n739) );
  NAND2_X1 U838 ( .A1(n745), .A2(n739), .ZN(n743) );
  INV_X1 U839 ( .A(n740), .ZN(n741) );
  OR2_X1 U840 ( .A1(n741), .A2(G286), .ZN(n742) );
  NAND2_X1 U841 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U843 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U844 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U845 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n753) );
  XNOR2_X1 U847 ( .A(n753), .B(KEYINPUT103), .ZN(n755) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  NOR2_X1 U849 ( .A1(n769), .A2(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  INV_X1 U851 ( .A(n774), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n1012), .A2(n767), .ZN(n757) );
  NOR2_X1 U853 ( .A1(n759), .A2(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U854 ( .A1(KEYINPUT33), .A2(n1011), .ZN(n760) );
  NOR2_X1 U855 ( .A1(n774), .A2(n760), .ZN(n761) );
  XNOR2_X1 U856 ( .A(n761), .B(KEYINPUT104), .ZN(n762) );
  NOR2_X1 U857 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U858 ( .A(n764), .B(KEYINPUT105), .ZN(n765) );
  NOR2_X1 U859 ( .A1(n1006), .A2(n765), .ZN(n778) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XNOR2_X1 U861 ( .A(KEYINPUT24), .B(n766), .ZN(n768) );
  NAND2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n776) );
  INV_X1 U863 ( .A(n769), .ZN(n772) );
  NOR2_X1 U864 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U865 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n812) );
  NAND2_X1 U870 ( .A1(G129), .A2(n889), .ZN(n780) );
  NAND2_X1 U871 ( .A1(G117), .A2(n890), .ZN(n779) );
  NAND2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n884), .A2(G105), .ZN(n781) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U876 ( .A(KEYINPUT93), .B(n784), .Z(n786) );
  NAND2_X1 U877 ( .A1(G141), .A2(n885), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n896) );
  AND2_X1 U879 ( .A1(n896), .A2(G1996), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G107), .A2(n890), .ZN(n788) );
  NAND2_X1 U881 ( .A1(G131), .A2(n885), .ZN(n787) );
  NAND2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U883 ( .A1(G119), .A2(n889), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G95), .A2(n884), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n878) );
  INV_X1 U887 ( .A(G1991), .ZN(n816) );
  NOR2_X1 U888 ( .A1(n878), .A2(n816), .ZN(n793) );
  NOR2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n950) );
  OR2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n827) );
  INV_X1 U892 ( .A(n827), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n950), .A2(n799), .ZN(n819) );
  XOR2_X1 U894 ( .A(KEYINPUT94), .B(n819), .Z(n810) );
  NAND2_X1 U895 ( .A1(n884), .A2(G104), .ZN(n801) );
  NAND2_X1 U896 ( .A1(G140), .A2(n885), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n802), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G128), .A2(n889), .ZN(n804) );
  NAND2_X1 U900 ( .A1(G116), .A2(n890), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U902 ( .A(n805), .B(KEYINPUT35), .Z(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U904 ( .A(KEYINPUT36), .B(n808), .Z(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT92), .B(n809), .Z(n879) );
  XNOR2_X1 U906 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NOR2_X1 U907 ( .A1(n879), .A2(n825), .ZN(n956) );
  NAND2_X1 U908 ( .A1(n827), .A2(n956), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n810), .A2(n822), .ZN(n811) );
  NOR2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n815) );
  XOR2_X1 U911 ( .A(G1986), .B(KEYINPUT91), .Z(n813) );
  XNOR2_X1 U912 ( .A(G290), .B(n813), .ZN(n1021) );
  NAND2_X1 U913 ( .A1(n1021), .A2(n827), .ZN(n814) );
  NAND2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n830) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n896), .ZN(n947) );
  AND2_X1 U916 ( .A1(n816), .A2(n878), .ZN(n952) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U918 ( .A1(n952), .A2(n817), .ZN(n818) );
  NOR2_X1 U919 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U920 ( .A1(n947), .A2(n820), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n824), .B(KEYINPUT106), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n879), .A2(n825), .ZN(n960) );
  NAND2_X1 U925 ( .A1(n826), .A2(n960), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U931 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G188) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(G325) );
  XNOR2_X1 U935 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(n838), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2474), .B(G1976), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1956), .B(G1981), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n841), .B(KEYINPUT110), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(G1971), .B(G1961), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1966), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2678), .Z(n851) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2090), .Z(n853) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U958 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U959 ( .A(G2096), .B(G2100), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U961 ( .A(G2078), .B(G2084), .Z(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U963 ( .A1(n889), .A2(G124), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G112), .A2(n890), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n884), .A2(G100), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G136), .A2(n885), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U970 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G127), .A2(n889), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G115), .A2(n890), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n869), .B(KEYINPUT47), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G103), .A2(n884), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G139), .A2(n885), .ZN(n872) );
  XNOR2_X1 U978 ( .A(KEYINPUT113), .B(n872), .ZN(n873) );
  NOR2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n962) );
  XNOR2_X1 U980 ( .A(G160), .B(n962), .ZN(n883) );
  XOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n876) );
  XNOR2_X1 U982 ( .A(G162), .B(KEYINPUT114), .ZN(n875) );
  XNOR2_X1 U983 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U984 ( .A(n953), .B(n877), .ZN(n881) );
  XNOR2_X1 U985 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U986 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U987 ( .A(n883), .B(n882), .ZN(n900) );
  NAND2_X1 U988 ( .A1(n884), .A2(G106), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G142), .A2(n885), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n888), .B(KEYINPUT45), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G130), .A2(n889), .ZN(n892) );
  NAND2_X1 U993 ( .A1(G118), .A2(n890), .ZN(n891) );
  NAND2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U995 ( .A(KEYINPUT112), .B(n893), .Z(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n897) );
  XOR2_X1 U997 ( .A(n897), .B(n896), .Z(n898) );
  XOR2_X1 U998 ( .A(G164), .B(n898), .Z(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n901), .ZN(G395) );
  XOR2_X1 U1001 ( .A(KEYINPUT115), .B(n902), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n903), .B(G171), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U1004 ( .A(G286), .B(n1019), .Z(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n908), .ZN(G397) );
  XOR2_X1 U1007 ( .A(G2451), .B(G2435), .Z(n910) );
  XNOR2_X1 U1008 ( .A(G2430), .B(G2454), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n916) );
  XOR2_X1 U1010 ( .A(G2427), .B(G2443), .Z(n912) );
  XNOR2_X1 U1011 ( .A(G1348), .B(G1341), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n914) );
  XOR2_X1 U1013 ( .A(G2446), .B(G2438), .Z(n913) );
  XNOR2_X1 U1014 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1015 ( .A(n916), .B(n915), .Z(n917) );
  NAND2_X1 U1016 ( .A1(G14), .A2(n917), .ZN(n923) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(n923), .ZN(G401) );
  XOR2_X1 U1025 ( .A(G2084), .B(G34), .Z(n924) );
  XNOR2_X1 U1026 ( .A(KEYINPUT54), .B(n924), .ZN(n941) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G35), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G26), .B(n925), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(G1996), .B(G32), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(G27), .B(n926), .ZN(n927) );
  NOR2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT118), .B(n933), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n934), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G25), .B(G1991), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(KEYINPUT53), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(KEYINPUT119), .ZN(n943) );
  XOR2_X1 U1043 ( .A(KEYINPUT55), .B(n943), .Z(n944) );
  NOR2_X1 U1044 ( .A1(G29), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n945), .B(KEYINPUT120), .ZN(n973) );
  INV_X1 U1046 ( .A(G29), .ZN(n971) );
  XOR2_X1 U1047 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1049 ( .A(KEYINPUT51), .B(n948), .Z(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G160), .B(G2084), .Z(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(KEYINPUT117), .B(n957), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n967) );
  XOR2_X1 U1058 ( .A(G2072), .B(n962), .Z(n964) );
  XOR2_X1 U1059 ( .A(G164), .B(G2078), .Z(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n965), .Z(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1063 ( .A(KEYINPUT52), .B(n968), .Z(n969) );
  NOR2_X1 U1064 ( .A1(KEYINPUT55), .A2(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1031) );
  XOR2_X1 U1067 ( .A(G16), .B(KEYINPUT124), .Z(n997) );
  XNOR2_X1 U1068 ( .A(G20), .B(n1008), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(G1981), .B(G6), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT59), .B(G1348), .Z(n978) );
  XNOR2_X1 U1074 ( .A(G4), .B(n978), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n981) );
  XNOR2_X1 U1077 ( .A(n982), .B(n981), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G21), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(G1961), .B(G5), .ZN(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G1986), .B(G24), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1085 ( .A(G1971), .B(KEYINPUT126), .Z(n989) );
  XNOR2_X1 U1086 ( .A(G22), .B(n989), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1088 ( .A(KEYINPUT58), .B(n992), .ZN(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(n995), .B(KEYINPUT61), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(G11), .A2(n998), .ZN(n1029) );
  XOR2_X1 U1093 ( .A(G16), .B(KEYINPUT56), .Z(n1027) );
  XNOR2_X1 U1094 ( .A(n1000), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(G1961), .B(KEYINPUT121), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(n1001), .B(G301), .ZN(n1002) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(n1004), .B(KEYINPUT122), .ZN(n1025) );
  XOR2_X1 U1099 ( .A(G1966), .B(G168), .Z(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1101 ( .A(KEYINPUT57), .B(n1007), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G303), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(KEYINPUT123), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(G1341), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(KEYINPUT127), .B(n1033), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

