//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NAND2_X1  g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT94), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  OAI22_X1  g008(.A1(new_n202), .A2(KEYINPUT15), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT95), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n209), .B(KEYINPUT93), .Z(new_n213));
  XNOR2_X1  g012(.A(new_n207), .B(KEYINPUT92), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n202), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(G8gat), .Z(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n217), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(KEYINPUT13), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G113gat), .B(G141gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G197gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT11), .B(G169gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n223), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n222), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n217), .A2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n225), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n227), .B(new_n234), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(KEYINPUT96), .ZN(new_n245));
  OR3_X1    g044(.A1(new_n240), .A2(KEYINPUT96), .A3(new_n241), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT97), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n245), .A2(KEYINPUT97), .A3(new_n243), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n247), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n227), .B1(new_n242), .B2(new_n243), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n233), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n257));
  INV_X1    g056(.A(G141gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G148gat), .ZN(new_n259));
  INV_X1    g058(.A(G148gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G141gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n259), .A2(new_n261), .B1(KEYINPUT2), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G155gat), .B(G162gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n262), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT78), .ZN(new_n267));
  INV_X1    g066(.A(G155gat), .ZN(new_n268));
  INV_X1    g067(.A(G162gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(KEYINPUT2), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n260), .A2(G141gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n258), .A2(G148gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n272), .A2(new_n276), .A3(KEYINPUT79), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT79), .B1(new_n272), .B2(new_n276), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n265), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(G211gat), .A2(G218gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(KEYINPUT22), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G211gat), .ZN(new_n284));
  INV_X1    g083(.A(G218gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT73), .A3(new_n281), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n287), .B(new_n280), .C1(KEYINPUT22), .C2(new_n282), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT29), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n279), .B1(KEYINPUT3), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT82), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n279), .B(new_n294), .C1(KEYINPUT3), .C2(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G228gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n265), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n303));
  INV_X1    g102(.A(new_n271), .ZN(new_n304));
  NOR3_X1   g103(.A1(KEYINPUT78), .A2(G155gat), .A3(G162gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n262), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n306), .B2(new_n263), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n272), .A2(new_n276), .A3(KEYINPUT79), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n289), .A2(new_n290), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n299), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n257), .B1(new_n296), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n299), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n300), .B1(new_n279), .B2(KEYINPUT3), .ZN(new_n316));
  INV_X1    g115(.A(new_n312), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n318), .A2(KEYINPUT83), .A3(new_n295), .A4(new_n293), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n286), .A2(new_n281), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n283), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n300), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n283), .A2(new_n322), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n310), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n279), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n299), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G22gat), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n332));
  INV_X1    g131(.A(G22gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n320), .A2(new_n333), .A3(new_n329), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n320), .B2(new_n329), .ZN(new_n336));
  AOI211_X1 g135(.A(G22gat), .B(new_n328), .C1(new_n314), .C2(new_n319), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT84), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT31), .B(G50gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n335), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G227gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n298), .ZN(new_n345));
  OR2_X1    g144(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(G183gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT65), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT24), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT65), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n346), .A2(new_n356), .A3(new_n347), .A4(new_n348), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT23), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n360), .A2(KEYINPUT25), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n360), .A2(new_n363), .A3(new_n362), .ZN(new_n367));
  OR2_X1    g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n355), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374));
  AND2_X1   g173(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G183gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT66), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n347), .A2(KEYINPUT27), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n374), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(new_n383), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT27), .B(G183gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT67), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n375), .A2(new_n376), .A3(new_n374), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n359), .A2(KEYINPUT26), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n351), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n363), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n359), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G113gat), .B(G120gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(KEYINPUT1), .ZN(new_n405));
  INV_X1    g204(.A(G134gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407));
  INV_X1    g206(.A(G127gat), .ZN(new_n408));
  INV_X1    g207(.A(G113gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G120gat), .ZN(new_n410));
  INV_X1    g209(.A(G120gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(G113gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n407), .B(new_n408), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n405), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n405), .B2(new_n413), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n373), .A2(new_n401), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n411), .A2(G113gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n409), .A2(G120gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n402), .B1(new_n420), .B2(new_n407), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT1), .B(G127gat), .C1(new_n418), .C2(new_n419), .ZN(new_n422));
  OAI21_X1  g221(.A(G134gat), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n358), .A2(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n399), .B1(new_n385), .B2(new_n392), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n345), .B1(new_n417), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT34), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT34), .B(new_n345), .C1(new_n417), .C2(new_n428), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT69), .ZN(new_n435));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT70), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n435), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n428), .A3(new_n345), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n439), .B(KEYINPUT32), .C1(new_n440), .C2(new_n438), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n433), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n433), .B1(new_n443), .B2(new_n444), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n336), .A2(new_n337), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n332), .A3(new_n341), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n343), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G226gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n298), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n426), .A2(new_n427), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(KEYINPUT29), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT75), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n457), .B(new_n453), .C1(new_n426), .C2(new_n427), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n379), .A2(new_n383), .A3(KEYINPUT67), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT67), .B1(new_n379), .B2(new_n383), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n377), .B(new_n381), .C1(new_n389), .C2(new_n380), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(new_n391), .B1(new_n463), .B2(new_n374), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n349), .A2(KEYINPUT65), .B1(new_n352), .B2(new_n354), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n364), .B1(new_n465), .B2(new_n357), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT25), .B1(new_n367), .B2(new_n369), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n464), .A2(new_n399), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n457), .B1(new_n468), .B2(new_n453), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n456), .B(new_n312), .C1(new_n459), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n453), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n301), .B1(new_n373), .B2(new_n401), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(new_n453), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n317), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n474), .A3(KEYINPUT76), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n458), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT76), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n312), .A4(new_n456), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G8gat), .B(G36gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n481), .B(new_n482), .Z(new_n483));
  AOI21_X1  g282(.A(KEYINPUT30), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT0), .ZN(new_n486));
  XNOR2_X1  g285(.A(G57gat), .B(G85gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  NAND2_X1  g287(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n309), .A2(new_n310), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n416), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n425), .A2(new_n309), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n425), .A2(new_n309), .A3(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n491), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n416), .A2(new_n279), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n492), .ZN(new_n500));
  INV_X1    g299(.A(new_n495), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n425), .B1(KEYINPUT3), .B2(new_n279), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(new_n490), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT4), .B1(new_n416), .B2(new_n279), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n425), .A2(new_n309), .A3(new_n493), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(KEYINPUT81), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n425), .A2(new_n309), .A3(new_n509), .A4(new_n493), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n505), .A2(new_n508), .A3(new_n498), .A4(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n488), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n511), .ZN(new_n514));
  INV_X1    g313(.A(new_n488), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n503), .A2(new_n511), .A3(new_n488), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n484), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n521));
  INV_X1    g320(.A(new_n483), .ZN(new_n522));
  AOI211_X1 g321(.A(new_n521), .B(new_n522), .C1(new_n475), .C2(new_n479), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n475), .A2(new_n522), .A3(new_n479), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n523), .A2(KEYINPUT77), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT77), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n480), .A2(KEYINPUT30), .A3(new_n483), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n475), .A2(new_n522), .A3(new_n479), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n520), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT35), .B1(new_n451), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n451), .C2(new_n530), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  AND4_X1   g334(.A1(new_n535), .A2(new_n514), .A3(KEYINPUT6), .A4(new_n515), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT86), .ZN(new_n539));
  AND4_X1   g338(.A1(new_n539), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT6), .B1(new_n514), .B2(new_n515), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n541), .B2(new_n518), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n443), .A2(new_n444), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n431), .A2(new_n432), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT71), .B1(new_n547), .B2(new_n445), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n433), .A2(new_n443), .A3(new_n444), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT71), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n484), .A2(new_n523), .A3(new_n524), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n543), .A2(new_n544), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n343), .A2(new_n450), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT89), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR4_X1   g355(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT84), .A4(new_n342), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n341), .B1(new_n449), .B2(new_n332), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n338), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n539), .A3(new_n518), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT35), .B1(new_n562), .B2(new_n538), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n446), .B2(new_n447), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n550), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n480), .A2(new_n483), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n521), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n528), .A3(new_n527), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT89), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n559), .A2(new_n563), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n533), .A2(new_n534), .A3(new_n556), .A4(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n574));
  AOI21_X1  g373(.A(new_n483), .B1(new_n480), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(new_n480), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT38), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n477), .A2(new_n317), .A3(new_n456), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n473), .B2(new_n312), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT38), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n575), .A2(new_n581), .B1(new_n483), .B2(new_n480), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n578), .A2(new_n562), .A3(new_n538), .A4(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n508), .A2(new_n491), .A3(new_n510), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n501), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n488), .B1(new_n586), .B2(KEYINPUT39), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT39), .B1(new_n500), .B2(new_n501), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n585), .B2(new_n501), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT85), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n587), .A2(new_n589), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n512), .B1(new_n593), .B2(KEYINPUT40), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n569), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n583), .A2(new_n595), .A3(new_n559), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT72), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n552), .B2(KEYINPUT36), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n448), .A2(KEYINPUT36), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n566), .A2(KEYINPUT72), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n530), .A2(new_n555), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n256), .B1(new_n573), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G71gat), .B(G78gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT98), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G57gat), .B(G64gat), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(KEYINPUT98), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n408), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n223), .B1(new_n612), .B2(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT99), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n268), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n619), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT7), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n632), .B1(new_n626), .B2(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G99gat), .B(G106gat), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n634), .B(KEYINPUT101), .ZN(new_n639));
  INV_X1    g438(.A(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(new_n612), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n612), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT102), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(KEYINPUT10), .A3(new_n612), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n643), .A2(new_n649), .A3(new_n644), .A4(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n643), .A2(new_n645), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n656), .A3(new_n660), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(G232gat), .A2(G233gat), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n642), .A2(new_n217), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n237), .A2(new_n638), .A3(new_n641), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(new_n239), .ZN(new_n668));
  XNOR2_X1  g467(.A(G190gat), .B(G218gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n665), .A2(KEYINPUT41), .ZN(new_n671));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n670), .B(new_n673), .Z(new_n674));
  NOR3_X1   g473(.A1(new_n625), .A2(new_n664), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n605), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n519), .A2(new_n513), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT103), .B(G1gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n569), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n682), .A2(G8gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n684), .B1(new_n690), .B2(new_n685), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g491(.A(G15gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n693), .A3(new_n552), .ZN(new_n694));
  INV_X1    g493(.A(new_n602), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n676), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(new_n693), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n676), .A2(new_n555), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND3_X1  g499(.A1(new_n556), .A2(new_n534), .A3(new_n572), .ZN(new_n701));
  INV_X1    g500(.A(new_n529), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n527), .A2(new_n526), .A3(new_n528), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n559), .A2(new_n704), .A3(new_n448), .A4(new_n520), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT90), .B1(new_n705), .B2(KEYINPUT35), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n604), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n674), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n664), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n625), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n256), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n674), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n710), .A2(KEYINPUT105), .A3(new_n713), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n677), .ZN(new_n720));
  INV_X1    g519(.A(new_n674), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n573), .B2(new_n604), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(new_n713), .ZN(new_n723));
  INV_X1    g522(.A(G29gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(new_n678), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n720), .A2(new_n726), .ZN(G1328gat));
  OAI21_X1  g526(.A(G36gat), .B1(new_n719), .B2(new_n553), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n712), .A2(G36gat), .A3(new_n721), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n605), .A2(new_n569), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1329gat));
  OAI21_X1  g531(.A(G43gat), .B1(new_n715), .B2(new_n602), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n566), .A2(G43gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n695), .A3(new_n718), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n737), .A2(new_n738), .A3(G43gat), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(G43gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n735), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n742), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g542(.A(G50gat), .B1(new_n715), .B2(new_n559), .ZN(new_n744));
  INV_X1    g543(.A(G50gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n723), .A2(new_n745), .A3(new_n555), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(KEYINPUT48), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n746), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n717), .A2(new_n555), .A3(new_n718), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(G50gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(G1331gat));
  NAND4_X1  g551(.A1(new_n256), .A2(new_n624), .A3(new_n721), .A4(new_n664), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n604), .B2(new_n573), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n678), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g555(.A(new_n553), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT108), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  INV_X1    g560(.A(G71gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n754), .A2(new_n762), .A3(new_n552), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n754), .A2(new_n695), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n762), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g565(.A1(new_n754), .A2(new_n555), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g567(.A1(new_n255), .A2(new_n711), .A3(new_n624), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n710), .A2(new_n714), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n710), .A2(KEYINPUT109), .A3(new_n714), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n677), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n255), .A2(new_n624), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n674), .A4(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n722), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n776), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n707), .A2(new_n674), .A3(new_n776), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n664), .A2(new_n626), .A3(new_n678), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n775), .B1(new_n785), .B2(new_n786), .ZN(G1336gat));
  OR2_X1    g586(.A1(new_n770), .A2(new_n553), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n627), .B1(new_n788), .B2(KEYINPUT112), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT112), .B2(new_n788), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n711), .A2(G92gat), .A3(new_n553), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n569), .A3(new_n773), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n781), .A2(new_n796), .A3(KEYINPUT51), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n781), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n795), .A2(G92gat), .B1(new_n799), .B2(new_n791), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n793), .B1(new_n794), .B2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n774), .B2(new_n602), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n711), .A2(G99gat), .A3(new_n566), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT113), .Z(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n785), .B2(new_n804), .ZN(G1338gat));
  NOR3_X1   g604(.A1(new_n711), .A2(G106gat), .A3(new_n559), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n784), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n784), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n710), .A2(new_n555), .A3(new_n714), .A4(new_n769), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n811), .B2(G106gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n806), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n797), .A2(new_n798), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n772), .A2(new_n555), .A3(new_n773), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(G106gat), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT115), .B(new_n813), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1339gat));
  NAND4_X1  g622(.A1(new_n647), .A2(new_n655), .A3(new_n648), .A4(new_n650), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n651), .A2(new_n826), .A3(new_n652), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n661), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n224), .A2(new_n226), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n241), .B2(new_n240), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n231), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n249), .B2(new_n250), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n661), .A4(new_n827), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n830), .A2(new_n834), .A3(new_n663), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n624), .B1(new_n836), .B2(new_n674), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n674), .B1(new_n834), .B2(new_n664), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n830), .A2(new_n663), .A3(new_n835), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n256), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n837), .A2(new_n840), .B1(new_n256), .B2(new_n675), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n677), .A3(new_n555), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(new_n448), .A3(new_n553), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n255), .A2(new_n409), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT116), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n570), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n256), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1340gat));
  NOR3_X1   g648(.A1(new_n847), .A2(new_n411), .A3(new_n711), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n843), .A2(new_n664), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n411), .ZN(G1341gat));
  NAND3_X1  g651(.A1(new_n843), .A2(new_n408), .A3(new_n624), .ZN(new_n853));
  OAI21_X1  g652(.A(G127gat), .B1(new_n847), .B2(new_n625), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1342gat));
  OAI21_X1  g654(.A(G134gat), .B1(new_n847), .B2(new_n721), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n721), .A2(new_n569), .ZN(new_n857));
  XOR2_X1   g656(.A(KEYINPUT68), .B(G134gat), .Z(new_n858));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n448), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(G1343gat));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n840), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n675), .A2(new_n256), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n555), .ZN(new_n869));
  XOR2_X1   g668(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n841), .B2(new_n559), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n602), .A2(new_n678), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n553), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n869), .A2(new_n871), .A3(new_n255), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G141gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n841), .A2(new_n559), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n256), .A2(G141gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n878), .A2(new_n553), .A3(new_n873), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n864), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n258), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n871), .A2(new_n875), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(KEYINPUT118), .A3(new_n255), .A4(new_n869), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n880), .A2(new_n864), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n882), .B(KEYINPUT119), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n884), .B2(new_n886), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n881), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n873), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n569), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n260), .A3(new_n664), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n867), .A2(new_n555), .A3(new_n870), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n867), .B2(new_n555), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n664), .B(new_n875), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n869), .A2(new_n871), .A3(new_n664), .A4(new_n875), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n902), .A2(new_n897), .A3(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n896), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT120), .B(new_n896), .C1(new_n901), .C2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n885), .A2(new_n869), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n624), .A2(G155gat), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT121), .Z(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G155gat), .B1(new_n895), .B2(new_n624), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT122), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n909), .B2(new_n721), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n857), .A2(new_n269), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n894), .B2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n553), .A2(new_n678), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n867), .A2(new_n552), .A3(new_n559), .A4(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(G169gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n256), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n867), .A2(new_n448), .A3(new_n559), .A4(new_n919), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n255), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n925), .B2(new_n921), .ZN(G1348gat));
  INV_X1    g725(.A(G176gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n927), .A3(new_n664), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n920), .B2(new_n711), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n920), .B2(new_n625), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n624), .A2(new_n462), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g733(.A(G190gat), .B1(new_n920), .B2(new_n721), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT61), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n377), .A3(new_n674), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1351gat));
  OR2_X1    g737(.A1(new_n898), .A2(new_n899), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n602), .A2(new_n919), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n942), .A2(new_n943), .A3(new_n256), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n878), .A2(new_n940), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n255), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n944), .A2(new_n946), .ZN(G1352gat));
  OAI21_X1  g746(.A(G204gat), .B1(new_n942), .B2(new_n711), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n711), .A2(G204gat), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n945), .A2(new_n949), .B1(KEYINPUT125), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n945), .A2(new_n284), .A3(new_n624), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n624), .A3(new_n941), .ZN(new_n958));
  AND4_X1   g757(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n284), .B1(KEYINPUT126), .B2(new_n960), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n958), .A2(new_n961), .B1(new_n957), .B2(KEYINPUT63), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n956), .B1(new_n959), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n942), .B2(new_n721), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n285), .A3(new_n674), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


