//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n468), .A2(G136), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT64), .A2(G114), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT64), .A2(G114), .ZN(new_n484));
  NOR3_X1   g059(.A1(new_n483), .A2(new_n484), .A3(new_n464), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n464), .C1(new_n480), .C2(new_n481), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n462), .A2(new_n490), .A3(G138), .A4(new_n464), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G651), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G651), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n494), .A2(new_n496), .A3(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G50), .ZN(new_n498));
  AND3_X1   g073(.A1(KEYINPUT65), .A2(KEYINPUT5), .A3(G543), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT5), .B1(KEYINPUT65), .B2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n494), .A2(new_n496), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G88), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n505));
  OAI21_X1  g080(.A(G62), .B1(new_n499), .B2(new_n500), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n505), .B1(new_n508), .B2(G651), .ZN(new_n509));
  AOI211_X1 g084(.A(KEYINPUT66), .B(new_n493), .C1(new_n506), .C2(new_n507), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n498), .B(new_n504), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT67), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT65), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT65), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT66), .B1(new_n518), .B2(new_n493), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n508), .A2(new_n505), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n521), .A2(new_n522), .A3(new_n498), .A4(new_n504), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n517), .A2(KEYINPUT68), .A3(G63), .A4(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n503), .A2(G89), .B1(new_n497), .B2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n497), .A2(G52), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n494), .A2(new_n496), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n517), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n493), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(G171));
  XOR2_X1   g117(.A(KEYINPUT69), .B(G43), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n497), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n537), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n493), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT70), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n497), .A2(G53), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n494), .A2(new_n496), .A3(G53), .A4(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n559), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n561), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(KEYINPUT73), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n568), .A2(KEYINPUT74), .A3(new_n493), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n568), .B2(new_n493), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n503), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(G299));
  OAI221_X1 g148(.A(new_n535), .B1(new_n537), .B2(new_n538), .C1(new_n540), .C2(new_n493), .ZN(G301));
  INV_X1    g149(.A(G166), .ZN(G303));
  AND2_X1   g150(.A1(new_n503), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(new_n497), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n497), .A2(G48), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n503), .A2(G86), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  OAI21_X1  g160(.A(G61), .B1(new_n499), .B2(new_n500), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n585), .B1(new_n588), .B2(G651), .ZN(new_n589));
  AOI211_X1 g164(.A(KEYINPUT75), .B(new_n493), .C1(new_n586), .C2(new_n587), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n583), .B(new_n584), .C1(new_n589), .C2(new_n590), .ZN(G305));
  XOR2_X1   g166(.A(KEYINPUT76), .B(G47), .Z(new_n592));
  AOI22_X1  g167(.A1(new_n503), .A2(G85), .B1(new_n497), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n593), .B(KEYINPUT77), .C1(new_n493), .C2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n497), .A2(new_n592), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n537), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n594), .A2(new_n493), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n595), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n537), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n503), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n497), .A2(KEYINPUT78), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n497), .A2(KEYINPUT78), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(G54), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(new_n493), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n608), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n603), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n603), .B1(new_n614), .B2(G868), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n569), .A2(new_n570), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n572), .B1(new_n563), .B2(new_n566), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n614), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n462), .A2(new_n469), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n474), .A2(G123), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT80), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n468), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT82), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT81), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n649), .B(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT83), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(KEYINPUT84), .ZN(new_n664));
  OAI21_X1  g239(.A(KEYINPUT17), .B1(new_n664), .B2(new_n658), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(new_n660), .Z(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n658), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(G2096), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(G2096), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT87), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n675), .A2(new_n678), .A3(new_n682), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n680), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(G166), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G16), .B2(G22), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G1971), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n694), .B(new_n697), .C1(G16), .C2(G22), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT32), .B(G1981), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n700), .A2(G23), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n581), .B2(new_n700), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(KEYINPUT33), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(KEYINPUT33), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G1976), .ZN(new_n714));
  INV_X1    g289(.A(G1976), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n711), .A2(new_n715), .A3(new_n712), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n699), .A2(new_n708), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n699), .A2(new_n717), .A3(new_n708), .A4(new_n719), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n700), .A2(G24), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n595), .A2(new_n601), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n700), .ZN(new_n727));
  MUX2_X1   g302(.A(new_n725), .B(new_n727), .S(KEYINPUT91), .Z(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G1986), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G25), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n474), .A2(G119), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT88), .ZN(new_n733));
  OR2_X1    g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n468), .A2(G131), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT90), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n731), .B1(new_n739), .B2(new_n730), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT35), .B(G1991), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G1986), .B2(new_n728), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n723), .A2(new_n724), .A3(new_n729), .A4(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n721), .A2(new_n729), .A3(new_n722), .A4(new_n745), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT36), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n730), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n730), .ZN(new_n752));
  MUX2_X1   g327(.A(new_n751), .B(new_n752), .S(KEYINPUT100), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(G171), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G5), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  NOR2_X1   g333(.A1(G164), .A2(new_n730), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G27), .B2(new_n730), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n757), .A2(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n763), .B1(new_n761), .B2(new_n760), .C1(G2090), .C2(new_n754), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n468), .A2(G139), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n469), .A2(G103), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT97), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n765), .B(new_n768), .C1(new_n770), .C2(new_n464), .ZN(new_n771));
  MUX2_X1   g346(.A(G33), .B(new_n771), .S(G29), .Z(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G2072), .Z(new_n773));
  XOR2_X1   g348(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n700), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n620), .B2(new_n700), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT102), .B(G1956), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n730), .A2(G32), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n468), .A2(G141), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n474), .A2(G129), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n469), .A2(G105), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n782), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT27), .B(G1996), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n773), .A2(new_n780), .A3(new_n781), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n700), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G168), .B2(new_n700), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G1966), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n730), .A2(G26), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n468), .A2(G140), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n474), .A2(G128), .ZN(new_n802));
  NOR2_X1   g377(.A1(G104), .A2(G2105), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n801), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n800), .B1(new_n805), .B2(G29), .ZN(new_n806));
  MUX2_X1   g381(.A(new_n800), .B(new_n806), .S(KEYINPUT28), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT95), .B(G2067), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n700), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n614), .B2(new_n700), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(G1348), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(G1348), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n809), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n549), .A2(new_n700), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n700), .B2(G19), .ZN(new_n816));
  INV_X1    g391(.A(G1341), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(KEYINPUT24), .A2(G34), .ZN(new_n819));
  NAND2_X1  g394(.A1(KEYINPUT24), .A2(G34), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n819), .A2(new_n730), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G160), .B2(new_n730), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G2084), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n639), .A2(new_n730), .ZN(new_n824));
  INV_X1    g399(.A(G28), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT30), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(KEYINPUT30), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(new_n827), .A3(new_n730), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n818), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT31), .B(G11), .Z(new_n830));
  OAI22_X1  g405(.A1(new_n816), .A2(new_n817), .B1(new_n757), .B2(new_n758), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n822), .A2(G2084), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT99), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n792), .A2(new_n794), .B1(new_n798), .B2(G1966), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n814), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NOR4_X1   g411(.A1(new_n764), .A2(new_n796), .A3(new_n799), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n750), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n748), .A2(KEYINPUT36), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n748), .B(new_n724), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(KEYINPUT36), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n841), .B2(KEYINPUT94), .ZN(G311));
  INV_X1    g417(.A(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n746), .A2(new_n749), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n845));
  OAI211_X1 g420(.A(KEYINPUT94), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n750), .A3(new_n837), .ZN(G150));
  AOI22_X1  g422(.A1(new_n503), .A2(G93), .B1(new_n497), .B2(G55), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(KEYINPUT103), .C1(new_n493), .C2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n497), .A2(G55), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n537), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n849), .A2(new_n493), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g431(.A(new_n544), .B1(new_n537), .B2(new_n545), .C1(new_n547), .C2(new_n493), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n850), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n854), .A2(new_n855), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n549), .A2(new_n859), .A3(KEYINPUT103), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n608), .A2(new_n611), .A3(new_n613), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n623), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  AOI21_X1  g442(.A(G860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n868), .B(new_n869), .C1(new_n867), .C2(new_n866), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT105), .ZN(new_n871));
  INV_X1    g446(.A(new_n859), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(G145));
  XNOR2_X1  g450(.A(new_n471), .B(new_n478), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n489), .A2(new_n491), .ZN(new_n877));
  OR2_X1    g452(.A1(KEYINPUT64), .A2(G114), .ZN(new_n878));
  NAND2_X1  g453(.A1(KEYINPUT64), .A2(G114), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(G2105), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n486), .ZN(new_n881));
  AOI22_X1  g456(.A1(G126), .A2(new_n474), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n805), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n876), .B(new_n884), .Z(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n468), .A2(G142), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n474), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n739), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n631), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n892), .A2(new_n631), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n886), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n893), .A3(new_n885), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n791), .B(KEYINPUT106), .Z(new_n900));
  MUX2_X1   g475(.A(new_n900), .B(new_n789), .S(new_n771), .Z(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(new_n639), .Z(new_n902));
  OR2_X1    g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n902), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g482(.A1(new_n872), .A2(G868), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n861), .B(new_n625), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n567), .A2(new_n863), .A3(new_n571), .A4(new_n572), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n910), .B2(new_n911), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT108), .B1(new_n620), .B2(new_n863), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n912), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n915), .B(new_n916), .C1(new_n909), .C2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n927));
  NAND2_X1  g502(.A1(G166), .A2(G290), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n581), .B(KEYINPUT109), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n726), .A2(new_n523), .A3(new_n512), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n933), .A2(new_n934), .A3(G305), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n929), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n702), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n927), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n926), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n908), .B1(new_n949), .B2(G868), .ZN(G295));
  AOI21_X1  g525(.A(new_n908), .B1(new_n949), .B2(G868), .ZN(G331));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  NAND4_X1  g527(.A1(G301), .A2(new_n531), .A3(new_n529), .A4(new_n532), .ZN(new_n953));
  NAND2_X1  g528(.A1(G286), .A2(G171), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n861), .A2(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n858), .A2(new_n860), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n924), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n937), .A2(new_n702), .A3(new_n932), .ZN(new_n960));
  OAI21_X1  g535(.A(G305), .B1(new_n933), .B2(new_n934), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n912), .B1(new_n956), .B2(new_n957), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n861), .B(new_n955), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n921), .B2(new_n923), .ZN(new_n965));
  INV_X1    g540(.A(new_n962), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n935), .A2(new_n938), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n967), .A3(new_n904), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n965), .A2(new_n966), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n939), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(KEYINPUT111), .A3(new_n912), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n962), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n922), .A2(new_n917), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n977), .A2(new_n958), .A3(new_n978), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n976), .A2(new_n979), .B1(new_n935), .B2(new_n938), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n972), .A2(KEYINPUT43), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n952), .B1(new_n970), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(new_n969), .A3(new_n980), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT44), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n982), .A2(new_n985), .A3(KEYINPUT112), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n970), .A2(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT44), .ZN(new_n989));
  AND4_X1   g564(.A1(new_n969), .A2(new_n980), .A3(new_n904), .A4(new_n963), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n969), .B1(new_n972), .B2(new_n967), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n952), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n986), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(KEYINPUT125), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT115), .B1(G164), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n877), .B2(new_n882), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT113), .B(G40), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n465), .A2(new_n470), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1966), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g583(.A(KEYINPUT119), .B(G1966), .C1(new_n1002), .C2(new_n1005), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1000), .B1(new_n883), .B2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT115), .B(G1384), .C1(new_n877), .C2(new_n882), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G2084), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n465), .A2(new_n470), .A3(new_n1003), .ZN(new_n1016));
  INV_X1    g591(.A(new_n999), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1008), .A2(new_n1009), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G168), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n1024), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT119), .B1(new_n1028), .B2(G1966), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1006), .A2(new_n996), .A3(new_n1007), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1019), .A3(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT51), .B(G8), .C1(new_n1031), .C2(G286), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT62), .B(new_n1025), .C1(new_n1027), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G2078), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1017), .A2(new_n998), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n999), .A2(KEYINPUT45), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1016), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1034), .B1(new_n1039), .B2(G2078), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1014), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n758), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1036), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT116), .B(G2090), .Z(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1014), .A2(new_n1016), .A3(new_n1018), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1039), .A2(new_n697), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1022), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(G166), .B2(new_n1022), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n512), .A2(new_n523), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G305), .A2(G1981), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT75), .B1(new_n1056), .B2(new_n493), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n588), .A2(new_n585), .A3(G651), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n583), .A4(new_n584), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1061), .A3(KEYINPUT49), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1055), .A2(new_n1061), .A3(new_n1067), .A4(KEYINPUT49), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n997), .A2(new_n1001), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1022), .B1(new_n1069), .B2(new_n1016), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1072));
  OAI221_X1 g647(.A(G8), .B1(new_n715), .B2(G288), .C1(new_n1072), .C2(new_n1004), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT52), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT117), .B(G1976), .Z(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1070), .B(new_n1076), .C1(new_n715), .C2(G288), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n997), .A2(KEYINPUT50), .A3(new_n1001), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n999), .A2(new_n1010), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1016), .A4(new_n1046), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1022), .B1(new_n1081), .B2(new_n1048), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1053), .ZN(new_n1083));
  NOR4_X1   g658(.A1(new_n1044), .A2(new_n1054), .A3(new_n1078), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n995), .B1(new_n1033), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1025), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1025), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT125), .A3(new_n1084), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1086), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1071), .A2(new_n715), .A3(new_n581), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1061), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1078), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1096), .A2(new_n1070), .B1(new_n1097), .B2(new_n1054), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1054), .A2(new_n1078), .A3(new_n1083), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1031), .A2(G8), .A3(G168), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT63), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT63), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1103));
  NOR4_X1   g678(.A1(new_n1100), .A2(new_n1103), .A3(new_n1054), .A4(new_n1078), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1098), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n563), .B2(new_n566), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g688(.A(G299), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1113), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(new_n620), .A3(new_n1111), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1079), .A2(new_n1080), .A3(new_n1016), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1039), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1117), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1118), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1127), .B(new_n1117), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1106), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1117), .A2(KEYINPUT123), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1114), .A2(new_n1116), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1121), .A2(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT61), .B(new_n1131), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1069), .A2(new_n1016), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(G2067), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1041), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1143), .A3(KEYINPUT60), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n614), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n863), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1148), .B2(new_n1144), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1140), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT58), .B(G1341), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1150), .A2(new_n1151), .B1(G1996), .B2(new_n1039), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n549), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT59), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1133), .A2(new_n1139), .A3(new_n1149), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1132), .A2(new_n863), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(new_n1146), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1042), .A2(new_n1040), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(G160), .B2(G40), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n465), .A2(new_n1162), .A3(G40), .A4(new_n470), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1035), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1161), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(G171), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(KEYINPUT54), .C1(G171), .C2(new_n1043), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1099), .A2(new_n1168), .ZN(new_n1169));
  OR3_X1    g744(.A1(new_n1160), .A2(G171), .A3(new_n1166), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT54), .B1(new_n1170), .B2(new_n1044), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1087), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1105), .B1(new_n1159), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1094), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n805), .B(G2067), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n791), .A2(G1996), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1175), .B(new_n1176), .C1(G1996), .C2(new_n789), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1016), .A2(new_n1017), .A3(new_n998), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT114), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1178), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n739), .A2(new_n742), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n739), .A2(new_n742), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(G290), .B(G1986), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1174), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT46), .ZN(new_n1190));
  OR3_X1    g765(.A1(new_n1178), .A2(new_n1190), .A3(G1996), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1182), .B1(new_n1175), .B2(new_n789), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1190), .B1(new_n1178), .B2(G1996), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT47), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1196));
  NOR2_X1   g771(.A1(G290), .A2(G1986), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1197), .A2(new_n1182), .A3(KEYINPUT48), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1181), .A2(new_n1199), .A3(new_n1185), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1182), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT48), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1196), .A2(new_n1198), .A3(new_n1200), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n805), .A2(G2067), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1205), .B1(new_n1208), .B2(new_n1182), .ZN(new_n1209));
  AOI211_X1 g784(.A(KEYINPUT126), .B(new_n1178), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1210));
  OAI211_X1 g785(.A(new_n1195), .B(new_n1204), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1189), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g788(.A(G401), .B1(new_n671), .B2(new_n672), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n983), .A2(new_n984), .ZN(new_n1216));
  NOR2_X1   g790(.A1(G229), .A2(new_n460), .ZN(new_n1217));
  NAND4_X1  g791(.A1(new_n906), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(G225));
  INV_X1    g792(.A(G225), .ZN(G308));
endmodule


