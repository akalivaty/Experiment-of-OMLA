

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n708), .A2(n707), .ZN(n712) );
  INV_X1 U554 ( .A(n735), .ZN(n704) );
  AND2_X1 U555 ( .A1(n542), .A2(n541), .ZN(n879) );
  BUF_X1 U556 ( .A(n880), .Z(n519) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n540), .Z(n880) );
  NAND2_X1 U558 ( .A1(n523), .A2(n988), .ZN(n759) );
  NAND2_X1 U559 ( .A1(n524), .A2(n522), .ZN(n806) );
  AND2_X1 U560 ( .A1(n804), .A2(n814), .ZN(n520) );
  AND2_X1 U561 ( .A1(n520), .A2(n805), .ZN(n521) );
  OR2_X1 U562 ( .A1(n770), .A2(n769), .ZN(n522) );
  OR2_X1 U563 ( .A1(n770), .A2(n757), .ZN(n523) );
  AND2_X1 U564 ( .A1(n766), .A2(n765), .ZN(n524) );
  XNOR2_X1 U565 ( .A(n705), .B(KEYINPUT26), .ZN(n706) );
  INV_X1 U566 ( .A(G168), .ZN(n693) );
  OR2_X1 U567 ( .A1(n770), .A2(G1966), .ZN(n688) );
  XNOR2_X1 U568 ( .A(n688), .B(KEYINPUT93), .ZN(n730) );
  NAND2_X1 U569 ( .A1(n791), .A2(n790), .ZN(n735) );
  INV_X1 U570 ( .A(KEYINPUT84), .ZN(n686) );
  OR2_X1 U571 ( .A1(n760), .A2(n759), .ZN(n766) );
  XNOR2_X1 U572 ( .A(n687), .B(n686), .ZN(n790) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n637) );
  NOR2_X1 U574 ( .A1(G651), .A2(n645), .ZN(n643) );
  NOR2_X1 U575 ( .A1(n542), .A2(n541), .ZN(n876) );
  NOR2_X1 U576 ( .A1(n547), .A2(n546), .ZN(G164) );
  XOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .Z(n645) );
  NAND2_X1 U578 ( .A1(G51), .A2(n643), .ZN(n527) );
  INV_X1 U579 ( .A(G651), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G543), .A2(n530), .ZN(n525) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n525), .Z(n649) );
  NAND2_X1 U582 ( .A1(G63), .A2(n649), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U584 ( .A(KEYINPUT6), .B(n528), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n637), .A2(G89), .ZN(n529) );
  XNOR2_X1 U586 ( .A(n529), .B(KEYINPUT4), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n645), .A2(n530), .ZN(n633) );
  NAND2_X1 U588 ( .A1(G76), .A2(n633), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U590 ( .A(n533), .B(KEYINPUT5), .Z(n534) );
  NOR2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U592 ( .A(KEYINPUT70), .B(n536), .Z(n537) );
  XNOR2_X1 U593 ( .A(KEYINPUT7), .B(n537), .ZN(G168) );
  AND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U595 ( .A1(G114), .A2(n875), .ZN(n539) );
  INV_X1 U596 ( .A(G2105), .ZN(n542) );
  XNOR2_X1 U597 ( .A(G2104), .B(KEYINPUT64), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G126), .A2(n876), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n547) );
  NOR2_X1 U600 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  NAND2_X1 U601 ( .A1(G138), .A2(n880), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G102), .A2(n879), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT83), .B(n545), .Z(n546) );
  NAND2_X1 U605 ( .A1(G91), .A2(n637), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G78), .A2(n633), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G53), .A2(n643), .ZN(n551) );
  NAND2_X1 U609 ( .A1(G65), .A2(n649), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U611 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U612 ( .A1(G85), .A2(n637), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G72), .A2(n633), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G47), .A2(n643), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G60), .A2(n649), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  OR2_X1 U618 ( .A1(n559), .A2(n558), .ZN(G290) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  NAND2_X1 U623 ( .A1(G52), .A2(n643), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G64), .A2(n649), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G90), .A2(n637), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G77), .A2(n633), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT65), .B(n564), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT9), .B(n565), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(G171) );
  NAND2_X1 U632 ( .A1(n649), .A2(G62), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT77), .B(n568), .Z(n570) );
  NAND2_X1 U634 ( .A1(n643), .A2(G50), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT78), .B(n571), .Z(n575) );
  NAND2_X1 U637 ( .A1(G88), .A2(n637), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G75), .A2(n633), .ZN(n572) );
  AND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(G303) );
  NAND2_X1 U641 ( .A1(n875), .A2(G113), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G101), .A2(n879), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT23), .B(n576), .Z(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n685) );
  NAND2_X1 U645 ( .A1(G137), .A2(n519), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G125), .A2(n876), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n683) );
  NOR2_X1 U648 ( .A1(n685), .A2(n683), .ZN(G160) );
  XOR2_X1 U649 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  XOR2_X1 U650 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n582) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U652 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U653 ( .A(KEYINPUT66), .B(n583), .ZN(G223) );
  XOR2_X1 U654 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n585) );
  INV_X1 U655 ( .A(G223), .ZN(n824) );
  NAND2_X1 U656 ( .A1(n824), .A2(G567), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n585), .B(n584), .ZN(G234) );
  NAND2_X1 U658 ( .A1(n637), .A2(G81), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G68), .A2(n633), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U662 ( .A(n589), .B(KEYINPUT13), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G43), .A2(n643), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n649), .A2(G56), .ZN(n592) );
  XOR2_X1 U666 ( .A(KEYINPUT14), .B(n592), .Z(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n970) );
  NAND2_X1 U668 ( .A1(n970), .A2(G860), .ZN(G153) );
  INV_X1 U669 ( .A(G171), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G54), .A2(n643), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G92), .A2(n637), .ZN(n596) );
  NAND2_X1 U673 ( .A1(G79), .A2(n633), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G66), .A2(n649), .ZN(n597) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(n597), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT15), .ZN(n979) );
  OR2_X1 U680 ( .A1(n979), .A2(G868), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U682 ( .A1(G868), .A2(G286), .ZN(n606) );
  INV_X1 U683 ( .A(G868), .ZN(n663) );
  NAND2_X1 U684 ( .A1(G299), .A2(n663), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(G297) );
  INV_X1 U686 ( .A(G860), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n607), .A2(G559), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n608), .A2(n979), .ZN(n609) );
  XNOR2_X1 U689 ( .A(n609), .B(KEYINPUT16), .ZN(n610) );
  XOR2_X1 U690 ( .A(KEYINPUT71), .B(n610), .Z(G148) );
  NAND2_X1 U691 ( .A1(n979), .A2(G868), .ZN(n611) );
  NOR2_X1 U692 ( .A1(G559), .A2(n611), .ZN(n613) );
  AND2_X1 U693 ( .A1(n663), .A2(n970), .ZN(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G111), .A2(n875), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G135), .A2(n519), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G123), .A2(n876), .ZN(n616) );
  XNOR2_X1 U699 ( .A(n616), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n879), .A2(G99), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n941) );
  XNOR2_X1 U703 ( .A(n941), .B(G2096), .ZN(n621) );
  XNOR2_X1 U704 ( .A(n621), .B(KEYINPUT72), .ZN(n623) );
  INV_X1 U705 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G93), .A2(n637), .ZN(n625) );
  NAND2_X1 U708 ( .A1(G80), .A2(n633), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G55), .A2(n643), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G67), .A2(n649), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U713 ( .A(KEYINPUT73), .B(n628), .Z(n629) );
  NOR2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n662) );
  NAND2_X1 U715 ( .A1(n979), .A2(G559), .ZN(n660) );
  XOR2_X1 U716 ( .A(n970), .B(n660), .Z(n631) );
  NOR2_X1 U717 ( .A1(G860), .A2(n631), .ZN(n632) );
  XNOR2_X1 U718 ( .A(n662), .B(n632), .ZN(G145) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(G73), .A2(n633), .ZN(n634) );
  XNOR2_X1 U721 ( .A(n634), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G48), .A2(n643), .ZN(n636) );
  NAND2_X1 U723 ( .A1(G61), .A2(n649), .ZN(n635) );
  NAND2_X1 U724 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n637), .A2(G86), .ZN(n638) );
  XOR2_X1 U726 ( .A(KEYINPUT76), .B(n638), .Z(n639) );
  NOR2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G49), .A2(n643), .ZN(n644) );
  XNOR2_X1 U730 ( .A(n644), .B(KEYINPUT74), .ZN(n651) );
  NAND2_X1 U731 ( .A1(G87), .A2(n645), .ZN(n647) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U736 ( .A(KEYINPUT75), .B(n652), .Z(G288) );
  XNOR2_X1 U737 ( .A(G290), .B(G305), .ZN(n658) );
  XNOR2_X1 U738 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U739 ( .A(G299), .B(n662), .ZN(n653) );
  XNOR2_X1 U740 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U741 ( .A(n970), .B(n655), .ZN(n656) );
  XNOR2_X1 U742 ( .A(n656), .B(G288), .ZN(n657) );
  XNOR2_X1 U743 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U744 ( .A(G166), .B(n659), .ZN(n896) );
  XNOR2_X1 U745 ( .A(n660), .B(n896), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n661), .A2(G868), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U749 ( .A(KEYINPUT80), .B(n666), .Z(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n667), .B(KEYINPUT81), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n668), .B(KEYINPUT20), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n669), .A2(G2090), .ZN(n670) );
  XNOR2_X1 U754 ( .A(n670), .B(KEYINPUT21), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n671), .B(KEYINPUT82), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U760 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G96), .A2(n675), .ZN(n829) );
  NAND2_X1 U762 ( .A1(n829), .A2(G2106), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U764 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U765 ( .A1(G108), .A2(n677), .ZN(n830) );
  NAND2_X1 U766 ( .A1(n830), .A2(G567), .ZN(n678) );
  NAND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n831) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U769 ( .A1(n831), .A2(n680), .ZN(n828) );
  NAND2_X1 U770 ( .A1(n828), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U772 ( .A1(G1971), .A2(G303), .ZN(n681) );
  NOR2_X1 U773 ( .A1(n756), .A2(n681), .ZN(n983) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n791) );
  INV_X1 U775 ( .A(G40), .ZN(n682) );
  OR2_X1 U776 ( .A1(n683), .A2(n682), .ZN(n684) );
  OR2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G8), .A2(n735), .ZN(n770) );
  INV_X1 U779 ( .A(KEYINPUT92), .ZN(n690) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n735), .ZN(n689) );
  XNOR2_X1 U781 ( .A(n690), .B(n689), .ZN(n731) );
  NAND2_X1 U782 ( .A1(G8), .A2(n731), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n730), .A2(n691), .ZN(n692) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT30), .ZN(n694) );
  AND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U786 ( .A(n695), .B(KEYINPUT97), .ZN(n699) );
  XOR2_X1 U787 ( .A(G2078), .B(KEYINPUT25), .Z(n929) );
  NOR2_X1 U788 ( .A1(n929), .A2(n735), .ZN(n697) );
  NOR2_X1 U789 ( .A1(n704), .A2(G1961), .ZN(n696) );
  NOR2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n726) );
  NAND2_X1 U791 ( .A1(n726), .A2(G301), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT31), .ZN(n742) );
  NOR2_X1 U794 ( .A1(G2067), .A2(n735), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n704), .A2(G1348), .ZN(n701) );
  NOR2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U797 ( .A1(G1341), .A2(n735), .ZN(n703) );
  XOR2_X1 U798 ( .A(KEYINPUT94), .B(n703), .Z(n708) );
  NAND2_X1 U799 ( .A1(n704), .A2(G1996), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n970), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n712), .A2(n979), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n711), .B(KEYINPUT95), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n979), .A2(n712), .ZN(n713) );
  NOR2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n720) );
  NAND2_X1 U806 ( .A1(n704), .A2(G2072), .ZN(n715) );
  XOR2_X1 U807 ( .A(KEYINPUT27), .B(n715), .Z(n717) );
  NAND2_X1 U808 ( .A1(G1956), .A2(n735), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G299), .A2(n721), .ZN(n718) );
  XNOR2_X1 U811 ( .A(n718), .B(KEYINPUT96), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U813 ( .A1(G299), .A2(n721), .ZN(n722) );
  XOR2_X1 U814 ( .A(KEYINPUT28), .B(n722), .Z(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U816 ( .A(n725), .B(KEYINPUT29), .ZN(n728) );
  OR2_X1 U817 ( .A1(G301), .A2(n726), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n741) );
  AND2_X1 U819 ( .A1(n742), .A2(n741), .ZN(n729) );
  NOR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n734) );
  INV_X1 U821 ( .A(n731), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n732), .A2(G8), .ZN(n733) );
  NAND2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n751) );
  INV_X1 U824 ( .A(G8), .ZN(n740) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n770), .ZN(n737) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n744) );
  AND2_X1 U830 ( .A1(n741), .A2(n744), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n748) );
  INV_X1 U832 ( .A(n744), .ZN(n746) );
  AND2_X1 U833 ( .A1(G286), .A2(G8), .ZN(n745) );
  OR2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U836 ( .A(n749), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n761) );
  NAND2_X1 U838 ( .A1(n983), .A2(n761), .ZN(n754) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U840 ( .A(n973), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n770), .A2(n752), .ZN(n753) );
  AND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n755), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  XOR2_X1 U845 ( .A(G1981), .B(KEYINPUT98), .Z(n758) );
  XNOR2_X1 U846 ( .A(G305), .B(n758), .ZN(n988) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n761), .A2(n763), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n764), .A2(n770), .ZN(n765) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XNOR2_X1 U852 ( .A(n767), .B(KEYINPUT91), .ZN(n768) );
  XNOR2_X1 U853 ( .A(KEYINPUT24), .B(n768), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G107), .A2(n875), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G131), .A2(n519), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U857 ( .A1(G95), .A2(n879), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G119), .A2(n876), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U861 ( .A(KEYINPUT86), .B(n777), .Z(n888) );
  AND2_X1 U862 ( .A1(G1991), .A2(n888), .ZN(n789) );
  NAND2_X1 U863 ( .A1(n879), .A2(G105), .ZN(n779) );
  XNOR2_X1 U864 ( .A(KEYINPUT88), .B(KEYINPUT38), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n779), .B(n778), .ZN(n786) );
  NAND2_X1 U866 ( .A1(G141), .A2(n519), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G129), .A2(n876), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G117), .A2(n875), .ZN(n782) );
  XNOR2_X1 U870 ( .A(KEYINPUT87), .B(n782), .ZN(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U873 ( .A(KEYINPUT89), .B(n787), .ZN(n872) );
  INV_X1 U874 ( .A(G1996), .ZN(n807) );
  NOR2_X1 U875 ( .A1(n872), .A2(n807), .ZN(n788) );
  NOR2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n945) );
  INV_X1 U877 ( .A(n790), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n819) );
  XOR2_X1 U879 ( .A(n819), .B(KEYINPUT90), .Z(n793) );
  NOR2_X1 U880 ( .A1(n945), .A2(n793), .ZN(n810) );
  INV_X1 U881 ( .A(n810), .ZN(n804) );
  XNOR2_X1 U882 ( .A(KEYINPUT37), .B(G2067), .ZN(n816) );
  NAND2_X1 U883 ( .A1(G104), .A2(n879), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G140), .A2(n519), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT34), .B(KEYINPUT85), .Z(n796) );
  XNOR2_X1 U887 ( .A(n797), .B(n796), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G116), .A2(n875), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G128), .A2(n876), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U891 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n803), .ZN(n892) );
  NOR2_X1 U894 ( .A1(n816), .A2(n892), .ZN(n950) );
  NAND2_X1 U895 ( .A1(n819), .A2(n950), .ZN(n814) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n972) );
  NAND2_X1 U897 ( .A1(n972), .A2(n819), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n521), .ZN(n822) );
  XOR2_X1 U899 ( .A(KEYINPUT39), .B(KEYINPUT99), .Z(n813) );
  AND2_X1 U900 ( .A1(n807), .A2(n872), .ZN(n947) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n888), .ZN(n942) );
  NOR2_X1 U903 ( .A1(n808), .A2(n942), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n947), .A2(n811), .ZN(n812) );
  XNOR2_X1 U906 ( .A(n813), .B(n812), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n892), .A2(n816), .ZN(n817) );
  XNOR2_X1 U909 ( .A(n817), .B(KEYINPUT100), .ZN(n960) );
  NAND2_X1 U910 ( .A1(n818), .A2(n960), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U913 ( .A(KEYINPUT40), .B(n823), .ZN(G329) );
  NAND2_X1 U914 ( .A1(n824), .A2(G2106), .ZN(n825) );
  XNOR2_X1 U915 ( .A(n825), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U917 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(G188) );
  XNOR2_X1 U920 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n831), .ZN(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(G1966), .Z(n833) );
  XNOR2_X1 U928 ( .A(G1996), .B(G1991), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U930 ( .A(n834), .B(KEYINPUT41), .Z(n836) );
  XNOR2_X1 U931 ( .A(G1961), .B(G1971), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U933 ( .A(G1976), .B(G1981), .Z(n838) );
  XNOR2_X1 U934 ( .A(G1986), .B(G1956), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U936 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT108), .B(G2474), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U940 ( .A(G2090), .B(KEYINPUT106), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n845), .B(G2678), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2100), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G227) );
  NAND2_X1 U949 ( .A1(G100), .A2(n879), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G136), .A2(n519), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n860) );
  NAND2_X1 U952 ( .A1(G112), .A2(n875), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n854), .B(KEYINPUT110), .ZN(n858) );
  XOR2_X1 U954 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n856) );
  NAND2_X1 U955 ( .A1(G124), .A2(n876), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U960 ( .A(n941), .B(KEYINPUT113), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n871) );
  NAND2_X1 U962 ( .A1(G115), .A2(n875), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G127), .A2(n876), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT47), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G139), .A2(n519), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n879), .A2(G103), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT112), .B(n868), .Z(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n953) );
  XOR2_X1 U971 ( .A(n871), .B(n953), .Z(n874) );
  XNOR2_X1 U972 ( .A(G164), .B(n872), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n894) );
  NAND2_X1 U974 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n886) );
  NAND2_X1 U977 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G142), .A2(n519), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(KEYINPUT45), .B(n883), .ZN(n884) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n884), .ZN(n885) );
  NOR2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U983 ( .A(n887), .B(G162), .Z(n890) );
  XNOR2_X1 U984 ( .A(G160), .B(n888), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U986 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U988 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U989 ( .A(G286), .B(n896), .ZN(n898) );
  XNOR2_X1 U990 ( .A(G171), .B(n979), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U992 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U993 ( .A(KEYINPUT103), .B(G2438), .Z(n901) );
  XNOR2_X1 U994 ( .A(G2443), .B(KEYINPUT102), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U996 ( .A(n902), .B(G2427), .Z(n904) );
  XNOR2_X1 U997 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U999 ( .A(G2451), .B(KEYINPUT101), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G2430), .B(G2454), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G2435), .B(G2446), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1005 ( .A1(n911), .A2(G14), .ZN(n917) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G34), .B(KEYINPUT118), .Z(n919) );
  XNOR2_X1 U1016 ( .A(G2084), .B(KEYINPUT54), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n919), .B(n918), .ZN(n937) );
  XNOR2_X1 U1018 ( .A(G2090), .B(G35), .ZN(n935) );
  XNOR2_X1 U1019 ( .A(G25), .B(G1991), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n920), .B(KEYINPUT115), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G1996), .B(G32), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(G28), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(G2072), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(G33), .B(n924), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n932) );
  XOR2_X1 U1029 ( .A(G27), .B(n929), .Z(n930) );
  XNOR2_X1 U1030 ( .A(KEYINPUT117), .B(n930), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT53), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT55), .B(n938), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(G29), .A2(n939), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(KEYINPUT119), .ZN(n968) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(KEYINPUT114), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n962) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT51), .B(n948), .Z(n952) );
  XOR2_X1 U1044 ( .A(G160), .B(G2084), .Z(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1047 ( .A(G2072), .B(n953), .Z(n955) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1050 ( .A(KEYINPUT50), .B(n956), .Z(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(n963), .B(KEYINPUT52), .ZN(n965) );
  INV_X1 U1055 ( .A(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(G29), .A2(n966), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n1024) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XOR2_X1 U1060 ( .A(G1956), .B(KEYINPUT121), .Z(n969) );
  XNOR2_X1 U1061 ( .A(G299), .B(n969), .ZN(n976) );
  XOR2_X1 U1062 ( .A(n970), .B(G1341), .Z(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n986) );
  XOR2_X1 U1068 ( .A(n979), .B(G1348), .Z(n981) );
  XOR2_X1 U1069 ( .A(G171), .B(G1961), .Z(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT120), .B(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(KEYINPUT122), .B(n987), .ZN(n992) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(KEYINPUT57), .B(n990), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n1021) );
  INV_X1 U1080 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n995), .B(G4), .ZN(n999) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G1956), .B(G20), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1087 ( .A(KEYINPUT123), .B(G1981), .Z(n1000) );
  XNOR2_X1 U1088 ( .A(G6), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(KEYINPUT124), .B(n1003), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1004), .B(KEYINPUT60), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G5), .B(G1961), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1016) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1012) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT125), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT126), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(G11), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(n1026), .B(KEYINPUT127), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

