//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n468), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(new_n465), .A2(new_n467), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(new_n475), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n481), .A2(new_n491), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT67), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n487), .A2(G126), .A3(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT69), .B1(new_n502), .B2(KEYINPUT68), .ZN(new_n503));
  OAI21_X1  g078(.A(G543), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(KEYINPUT69), .B(G543), .C1(new_n502), .C2(KEYINPUT68), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(G62), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n505), .A2(G88), .A3(new_n506), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(G50), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(G166));
  AND2_X1   g089(.A1(new_n510), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G51), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n505), .A2(G89), .A3(new_n506), .A4(new_n510), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n505), .A2(G63), .A3(G651), .A4(new_n506), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n516), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(G286));
  INV_X1    g096(.A(G286), .ZN(G168));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n523), .B2(KEYINPUT5), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n506), .B(new_n510), .C1(new_n525), .C2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n510), .A2(G543), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n505), .A2(G64), .A3(new_n506), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n501), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  OAI211_X1 g111(.A(G56), .B(new_n506), .C1(new_n525), .C2(new_n527), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n537), .A2(KEYINPUT70), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT70), .B1(new_n537), .B2(new_n538), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n505), .A2(G81), .A3(new_n506), .A4(new_n510), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n510), .A2(G43), .A3(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT71), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(KEYINPUT71), .A3(new_n543), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n541), .A2(G651), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n505), .A2(new_n556), .A3(new_n506), .A4(new_n510), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n559), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n505), .A2(G65), .A3(new_n506), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n501), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n558), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  AND2_X1   g143(.A1(new_n511), .A2(new_n512), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n507), .A2(new_n508), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(new_n501), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(G166), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G303));
  NAND2_X1  g150(.A1(new_n505), .A2(new_n506), .ZN(new_n576));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n501), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n555), .A2(new_n557), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT75), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(new_n583), .ZN(G288));
  NAND3_X1  g159(.A1(new_n505), .A2(G61), .A3(new_n506), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT76), .B1(new_n531), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n510), .A2(new_n591), .A3(G48), .A4(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n555), .B2(new_n557), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  NAND3_X1  g173(.A1(new_n505), .A2(G60), .A3(new_n506), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT77), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n599), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(G651), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n528), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G47), .B2(new_n515), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT78), .B1(G171), .B2(new_n610), .ZN(new_n611));
  OR3_X1    g186(.A1(G171), .A2(KEYINPUT78), .A3(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n579), .A2(G92), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n576), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n579), .A2(new_n619), .A3(G92), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n614), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n611), .B(new_n612), .C1(new_n622), .C2(G868), .ZN(G284));
  OAI211_X1 g198(.A(new_n611), .B(new_n612), .C1(new_n622), .C2(G868), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n566), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n566), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NOR3_X1   g204(.A1(new_n539), .A2(new_n540), .A3(new_n501), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n542), .A2(KEYINPUT71), .A3(new_n543), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(new_n544), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n610), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n622), .A2(new_n628), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT79), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n633), .B1(new_n635), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n479), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n481), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT81), .B(KEYINPUT82), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT16), .B(G2443), .Z(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n663), .A2(G14), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT17), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n672), .C2(new_n668), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT19), .Z(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(KEYINPUT84), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g262(.A(new_n683), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n680), .A2(new_n681), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT83), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1986), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1991), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n694), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G25), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n479), .A2(G119), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G131), .ZN(new_n703));
  OR2_X1    g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT35), .B(G1991), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  AND2_X1   g285(.A1(new_n605), .A2(new_n608), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n712), .B2(G24), .ZN(new_n714));
  INV_X1    g289(.A(G1986), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n712), .A2(G23), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G288), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT33), .Z(new_n719));
  INV_X1    g294(.A(G1976), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n718), .B(KEYINPUT33), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1976), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n712), .A2(G6), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n597), .B2(new_n712), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT32), .B(G1981), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n725), .A2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G22), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT85), .B1(new_n730), .B2(G16), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n730), .A2(KEYINPUT85), .A3(G16), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n731), .B(new_n732), .C1(G166), .C2(new_n712), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G1971), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n728), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n733), .A2(G1971), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n721), .A2(new_n723), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n716), .B1(new_n737), .B2(KEYINPUT34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n714), .A2(new_n715), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n738), .B(new_n739), .C1(KEYINPUT34), .C2(new_n737), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT36), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G11), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT90), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n479), .A2(G129), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n481), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G29), .B2(G32), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2072), .ZN(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  INV_X1    g332(.A(G127), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n468), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n759), .A2(G2105), .B1(new_n481), .B2(G139), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G29), .B2(G33), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n755), .B1(new_n756), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n756), .B2(new_n766), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n642), .A2(new_n700), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT30), .B(G28), .Z(new_n770));
  OAI221_X1 g345(.A(new_n769), .B1(G29), .B2(new_n770), .C1(new_n753), .C2(new_n754), .ZN(new_n771));
  INV_X1    g346(.A(G2078), .ZN(new_n772));
  NOR2_X1   g347(.A1(G164), .A2(new_n700), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G27), .B2(new_n700), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NOR2_X1   g351(.A1(KEYINPUT24), .A2(G34), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n700), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n780), .B(new_n781), .C1(new_n477), .C2(new_n700), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n742), .A2(new_n768), .A3(new_n775), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT89), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n700), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT87), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n479), .A2(G128), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n481), .A2(G140), .ZN(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n700), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n774), .B2(new_n772), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n712), .A2(G21), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G168), .B2(new_n712), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1966), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G171), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G5), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n785), .A2(new_n787), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT92), .B(KEYINPUT23), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n712), .A2(G20), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G299), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1956), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n807), .B2(new_n806), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n700), .A2(G35), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G162), .B2(new_n700), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT29), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2090), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n712), .A2(G4), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n622), .B2(new_n712), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1348), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n809), .A2(new_n817), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n712), .A2(G19), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n547), .B2(new_n712), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT86), .B(G1341), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n741), .A2(new_n825), .A3(new_n829), .ZN(G311));
  NAND3_X1  g405(.A1(new_n741), .A2(new_n825), .A3(new_n829), .ZN(G150));
  OAI211_X1 g406(.A(G67), .B(new_n506), .C1(new_n525), .C2(new_n527), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT95), .B1(new_n834), .B2(G651), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n528), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G55), .B2(new_n515), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(KEYINPUT95), .A3(G651), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n622), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n547), .A2(new_n841), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n847));
  AOI211_X1 g422(.A(new_n847), .B(new_n501), .C1(new_n832), .C2(new_n833), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n835), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(new_n839), .C1(new_n630), .C2(new_n632), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n853), .B2(KEYINPUT96), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(KEYINPUT96), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n843), .B1(new_n855), .B2(new_n856), .ZN(G145));
  INV_X1    g432(.A(new_n751), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n497), .B1(new_n490), .B2(new_n492), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n795), .A3(new_n496), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n795), .B1(new_n859), .B2(new_n496), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(new_n764), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n499), .A2(new_n796), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n763), .B1(new_n864), .B2(new_n860), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n858), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n764), .B1(new_n861), .B2(new_n862), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n763), .A3(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n751), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n479), .A2(G130), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n481), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(new_n645), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n706), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n866), .A2(new_n877), .A3(new_n869), .ZN(new_n880));
  XNOR2_X1  g455(.A(G160), .B(new_n642), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n485), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT98), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT97), .ZN(new_n889));
  INV_X1    g464(.A(new_n882), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n889), .B(new_n890), .C1(KEYINPUT97), .C2(new_n879), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT99), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n887), .A2(new_n894), .A3(new_n891), .A4(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n841), .A2(new_n610), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n635), .B(new_n851), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n621), .A2(G299), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n619), .B1(new_n579), .B2(G92), .ZN(new_n901));
  INV_X1    g476(.A(G92), .ZN(new_n902));
  AOI211_X1 g477(.A(KEYINPUT10), .B(new_n902), .C1(new_n555), .C2(new_n557), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n566), .A3(new_n618), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n900), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n900), .B2(new_n905), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n899), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(G166), .B1(new_n594), .B2(new_n596), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n579), .A2(G86), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n587), .A2(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n571), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G87), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n555), .B2(new_n557), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n924), .A2(new_n582), .A3(new_n578), .ZN(new_n925));
  NOR2_X1   g500(.A1(G290), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G290), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT101), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n922), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n916), .A2(new_n919), .ZN(new_n931));
  INV_X1    g506(.A(new_n928), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n931), .B(KEYINPUT101), .C1(new_n932), .C2(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(new_n934), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n915), .B(new_n940), .Z(new_n941));
  OAI21_X1  g516(.A(new_n898), .B1(new_n941), .B2(new_n610), .ZN(G295));
  OAI21_X1  g517(.A(new_n898), .B1(new_n941), .B2(new_n610), .ZN(G331));
  AOI21_X1  g518(.A(new_n566), .B1(new_n904), .B2(new_n618), .ZN(new_n944));
  AND4_X1   g519(.A1(new_n566), .A2(new_n614), .A3(new_n618), .A4(new_n620), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(G168), .B1(new_n535), .B2(new_n532), .ZN(new_n947));
  NAND2_X1  g522(.A1(G171), .A2(G286), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n846), .A2(new_n850), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n846), .B2(new_n850), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n846), .A2(new_n850), .A3(new_n949), .ZN(new_n955));
  INV_X1    g530(.A(new_n951), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n955), .B(new_n956), .C1(new_n909), .C2(new_n912), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n946), .B(KEYINPUT105), .C1(new_n950), .C2(new_n951), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n934), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n930), .A2(new_n933), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(new_n957), .A3(new_n962), .A4(new_n958), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n960), .A2(new_n961), .A3(new_n888), .A4(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n963), .A2(new_n888), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n967), .A2(KEYINPUT107), .A3(new_n961), .A4(new_n960), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n906), .B1(new_n956), .B2(new_n955), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n906), .A2(new_n908), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n900), .A2(new_n905), .A3(new_n910), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n956), .A3(new_n955), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n950), .A2(new_n951), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(KEYINPUT106), .A3(new_n971), .A4(new_n970), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n962), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n963), .A2(new_n888), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n966), .A2(new_n968), .A3(KEYINPUT44), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n973), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n952), .A3(new_n976), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n934), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n967), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n982), .B1(new_n986), .B2(KEYINPUT43), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n966), .A4(new_n968), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n981), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n961), .B1(new_n967), .B2(new_n960), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n995), .ZN(G397));
  AOI21_X1  g571(.A(G1384), .B1(new_n859), .B2(new_n496), .ZN(new_n997));
  NAND2_X1  g572(.A1(G160), .A2(G40), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n997), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT110), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n795), .B(new_n798), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n858), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1996), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT109), .Z(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(KEYINPUT46), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(KEYINPUT46), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1006), .A2(new_n858), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1001), .B1(new_n1004), .B2(new_n751), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1013));
  NOR4_X1   g588(.A1(new_n1011), .A2(new_n709), .A3(new_n706), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n795), .A2(G2067), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1000), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n706), .B(new_n709), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1013), .B(new_n1011), .C1(new_n1000), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G290), .A2(G1986), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n999), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1010), .A2(new_n1016), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1966), .ZN(new_n1024));
  OAI211_X1 g599(.A(G40), .B(G160), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1026), .B(G1384), .C1(new_n859), .C2(new_n496), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n499), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n997), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n477), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n783), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G286), .A2(G8), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT123), .B1(G286), .B2(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(KEYINPUT51), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(G8), .A3(G286), .ZN(new_n1044));
  OAI211_X1 g619(.A(G8), .B(new_n1041), .C1(new_n1037), .C2(G286), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT62), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1049));
  INV_X1    g624(.A(G2090), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1031), .A2(new_n1033), .A3(new_n1050), .A4(new_n1035), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(G303), .B2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1053), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1055), .B(new_n1056), .C1(new_n572), .C2(new_n574), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(G8), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n997), .B2(new_n1035), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G288), .A2(new_n720), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(new_n1061), .C1(new_n1062), .C2(KEYINPUT113), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(KEYINPUT113), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1060), .A2(KEYINPUT113), .A3(new_n720), .A4(G288), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1067), .B(new_n1066), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1052), .A2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1058), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n597), .A2(new_n696), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n528), .A2(new_n595), .ZN(new_n1076));
  OAI21_X1  g651(.A(G1981), .B1(new_n594), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(KEYINPUT115), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1081), .B(KEYINPUT49), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1078), .B(new_n1060), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  AND4_X1   g658(.A1(new_n1059), .A2(new_n1071), .A3(new_n1074), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1034), .B1(new_n1030), .B2(new_n1026), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n997), .A2(KEYINPUT45), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n772), .A3(G160), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1031), .A2(new_n1035), .A3(new_n1033), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1087), .A2(new_n1088), .B1(new_n807), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1027), .A2(new_n1088), .A3(G2078), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(G160), .A3(new_n1085), .ZN(new_n1092));
  AOI21_X1  g667(.A(G301), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1043), .A2(new_n1094), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1047), .A2(new_n1084), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1037), .A2(new_n1097), .A3(G8), .A4(G168), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1059), .ZN(new_n1099));
  AND4_X1   g674(.A1(new_n1074), .A2(new_n1099), .A3(new_n1083), .A4(new_n1071), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1060), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1083), .A2(new_n720), .A3(new_n925), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1075), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1072), .A2(KEYINPUT116), .A3(new_n1073), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1038), .A2(G286), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1052), .B(G8), .C1(new_n1107), .C2(new_n1058), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1071), .A2(new_n1083), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT63), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1096), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1113), .A2(new_n1114), .B1(new_n1089), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n566), .B1(KEYINPUT117), .B2(KEYINPUT57), .ZN(new_n1117));
  NOR2_X1   g692(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1089), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n499), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n997), .A2(KEYINPUT118), .A3(new_n1035), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n798), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n622), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1119), .B2(new_n1116), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n547), .A2(KEYINPUT121), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1025), .A2(G1996), .A3(new_n1027), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(G1341), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT120), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT118), .B1(new_n997), .B2(new_n1035), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1085), .A2(new_n1004), .A3(G160), .A4(new_n1086), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1131), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1146), .B(new_n1131), .C1(new_n1137), .C2(new_n1143), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1128), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n621), .B1(new_n1149), .B2(KEYINPUT60), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1128), .A2(new_n1151), .A3(new_n622), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1150), .A2(new_n1152), .B1(KEYINPUT60), .B2(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1130), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1155), .A2(new_n1129), .A3(new_n1156), .A4(KEYINPUT61), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1120), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n470), .A2(KEYINPUT124), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n470), .A2(KEYINPUT124), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n475), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1085), .A2(KEYINPUT125), .A3(new_n476), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n1166));
  OAI211_X1 g741(.A(G40), .B(new_n476), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n1163), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(new_n1091), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1090), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(G171), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1160), .B1(new_n1171), .B2(new_n1093), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1155), .A2(KEYINPUT61), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1172), .A2(new_n1084), .A3(new_n1173), .A4(new_n1046), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1090), .A2(new_n1169), .A3(KEYINPUT126), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(G171), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1090), .A2(G301), .A3(new_n1092), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1178), .A2(KEYINPUT54), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1112), .B1(new_n1159), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n711), .A2(new_n715), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n999), .B1(new_n1183), .B2(new_n1019), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1018), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT111), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1018), .A2(KEYINPUT111), .A3(new_n1184), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1023), .B1(new_n1182), .B2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g765(.A(G401), .B1(new_n893), .B2(new_n895), .ZN(new_n1192));
  NOR3_X1   g766(.A1(G229), .A2(new_n461), .A3(G227), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n993), .A2(new_n1192), .A3(new_n1193), .ZN(G308));
  NAND3_X1  g768(.A1(new_n993), .A2(new_n1192), .A3(new_n1193), .ZN(G225));
endmodule


