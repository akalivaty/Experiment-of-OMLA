//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT67), .Z(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(G126), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n464), .B2(new_n465), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n464), .B2(new_n465), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n497), .C1(new_n465), .C2(new_n464), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT69), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n500), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT70), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(new_n506), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n508), .B2(new_n500), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(G651), .B1(G50), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n520), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT7), .Z(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n527), .B2(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n513), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n513), .A2(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n506), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G651), .B1(G52), .B2(new_n520), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n513), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n506), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(G43), .B2(new_n520), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n506), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n507), .A2(new_n512), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n520), .A2(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(KEYINPUT73), .B2(KEYINPUT9), .ZN(new_n563));
  AND2_X1   g138(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n564));
  NOR2_X1   g139(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n520), .B(G53), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n563), .A2(KEYINPUT74), .A3(new_n566), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n561), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n522), .A2(KEYINPUT75), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n514), .A2(new_n574), .A3(new_n521), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(G303));
  OR2_X1    g151(.A1(new_n510), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n520), .B2(G49), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n559), .B2(new_n579), .ZN(G288));
  AND3_X1   g155(.A1(new_n507), .A2(G86), .A3(new_n512), .ZN(new_n581));
  OAI21_X1  g156(.A(G61), .B1(new_n504), .B2(new_n505), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n520), .A2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n520), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G651), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n590), .B1(new_n591), .B2(new_n592), .C1(new_n559), .C2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n520), .A2(G54), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n591), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n507), .A2(G92), .A3(new_n512), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(KEYINPUT10), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT76), .Z(new_n604));
  AOI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(new_n595), .ZN(G284));
  AOI21_X1  g180(.A(new_n596), .B1(new_n604), .B2(new_n595), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n571), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(G868), .B2(new_n571), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n604), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n477), .A2(G135), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n463), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n616), .B1(new_n617), .B2(new_n618), .C1(new_n619), .C2(new_n483), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n482), .A2(new_n471), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT77), .ZN(new_n627));
  AOI211_X1 g202(.A(new_n621), .B(new_n627), .C1(new_n625), .C2(new_n624), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT79), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n645), .B1(new_n647), .B2(KEYINPUT80), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(KEYINPUT80), .B2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2084), .B(G2090), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n647), .B(KEYINPUT17), .Z(new_n651));
  INV_X1    g226(.A(new_n645), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n645), .A2(new_n650), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n625), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT81), .B(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(KEYINPUT82), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(G229));
  NAND2_X1  g261(.A1(new_n482), .A2(G127), .ZN(new_n687));
  INV_X1    g262(.A(G115), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n470), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n463), .B1(new_n689), .B2(KEYINPUT89), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(KEYINPUT89), .B2(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT25), .Z(new_n693));
  AOI21_X1  g268(.A(KEYINPUT88), .B1(new_n477), .B2(G139), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n477), .A2(KEYINPUT88), .A3(G139), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n691), .B(new_n693), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  MUX2_X1   g271(.A(G33), .B(new_n696), .S(G29), .Z(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G2072), .Z(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G21), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G168), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G1966), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT29), .Z(new_n707));
  INV_X1    g282(.A(G2090), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n707), .A2(new_n708), .B1(new_n701), .B2(G1966), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n698), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n699), .A2(G4), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n604), .B2(new_n699), .ZN(new_n712));
  INV_X1    g287(.A(G1348), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n704), .A2(G32), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  INV_X1    g292(.A(G129), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n483), .B2(new_n718), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT90), .Z(new_n723));
  OAI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(new_n704), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT27), .B(G1996), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n548), .A2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G16), .B2(G19), .ZN(new_n728));
  INV_X1    g303(.A(G1341), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  NOR2_X1   g305(.A1(G5), .A2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT92), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G301), .B2(new_n699), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n730), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(new_n729), .C2(new_n728), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n737), .A2(new_n704), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n704), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n704), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n740), .B1(new_n704), .B2(new_n620), .C1(new_n742), .C2(G2078), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n704), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n704), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2084), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n704), .A2(G26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT87), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G116), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT86), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n477), .A2(G140), .ZN(new_n758));
  INV_X1    g333(.A(G128), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n483), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n704), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n762), .A2(G2067), .B1(G2078), .B2(new_n742), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n750), .B(new_n763), .C1(G2067), .C2(new_n762), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n726), .A2(new_n736), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n710), .A2(new_n714), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n699), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n708), .B2(new_n707), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n699), .A2(G22), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n699), .ZN(new_n776));
  INV_X1    g351(.A(G1971), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G6), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n588), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G23), .B(G288), .S(G16), .Z(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n778), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n704), .A2(G25), .ZN(new_n789));
  INV_X1    g364(.A(new_n483), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G119), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT84), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G107), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G131), .B2(new_n477), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(new_n704), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  XOR2_X1   g376(.A(new_n800), .B(new_n801), .Z(new_n802));
  MUX2_X1   g377(.A(G24), .B(G290), .S(G16), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1986), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n788), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(KEYINPUT85), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT85), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n788), .B2(new_n805), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n787), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT36), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(new_n787), .C1(new_n807), .C2(new_n809), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n774), .B1(new_n811), .B2(new_n813), .ZN(G311));
  XNOR2_X1  g389(.A(new_n806), .B(KEYINPUT85), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n812), .B1(new_n815), .B2(new_n787), .ZN(new_n816));
  INV_X1    g391(.A(new_n813), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n773), .B1(new_n816), .B2(new_n817), .ZN(G150));
  XOR2_X1   g393(.A(KEYINPUT95), .B(G93), .Z(new_n819));
  NOR2_X1   g394(.A1(new_n559), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n520), .A2(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n591), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n604), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n824), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n542), .A2(new_n832), .A3(new_n546), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n542), .B2(new_n546), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n837), .A2(new_n824), .A3(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n830), .B(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n825), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n827), .B1(new_n841), .B2(new_n842), .ZN(G145));
  NAND2_X1  g418(.A1(new_n496), .A2(new_n498), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n489), .B1(new_n475), .B2(new_n476), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n463), .A2(G114), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n845), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT97), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n844), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n761), .B(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n790), .A2(G130), .B1(G142), .B2(new_n477), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  INV_X1    g430(.A(G118), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n855), .A2(KEYINPUT98), .B1(new_n856), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(KEYINPUT98), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n853), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n798), .B(new_n623), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n722), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n696), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n723), .B2(new_n696), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n620), .B(G160), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G162), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n870), .A3(new_n867), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g451(.A1(new_n831), .A2(new_n595), .ZN(new_n877));
  XNOR2_X1  g452(.A(G290), .B(G288), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT101), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n522), .B(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(G305), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n522), .B(KEYINPUT100), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n588), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n879), .B(new_n880), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n588), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(G305), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT101), .A4(new_n878), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n890), .B2(KEYINPUT102), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n612), .A2(new_n839), .ZN(new_n897));
  INV_X1    g472(.A(new_n839), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n604), .A2(new_n610), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n603), .A2(new_n571), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n603), .A2(new_n571), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT99), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(new_n903), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(KEYINPUT41), .A3(new_n901), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n897), .A2(new_n899), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n912));
  INV_X1    g487(.A(new_n899), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n898), .B1(new_n604), .B2(new_n610), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n912), .B(new_n904), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n896), .A2(new_n906), .A3(new_n911), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n911), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n912), .B1(new_n900), .B2(new_n904), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n891), .B(new_n895), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n877), .B1(new_n920), .B2(new_n595), .ZN(G295));
  OAI21_X1  g496(.A(new_n877), .B1(new_n920), .B2(new_n595), .ZN(G331));
  XOR2_X1   g497(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(G286), .A2(G301), .ZN(new_n925));
  NAND2_X1  g500(.A1(G168), .A2(G171), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n836), .A2(new_n838), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n836), .A2(new_n838), .B1(new_n926), .B2(new_n925), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n908), .B(new_n910), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n839), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n904), .A3(new_n927), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n927), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n908), .A4(new_n910), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n938), .B2(new_n892), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n931), .A2(new_n890), .A3(new_n934), .A4(new_n937), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n924), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n930), .A2(new_n934), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(new_n892), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n943), .A2(new_n940), .A3(new_n924), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n923), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n892), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n924), .A3(new_n873), .A4(new_n940), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n940), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n943), .B2(new_n940), .ZN(new_n951));
  OAI211_X1 g526(.A(KEYINPUT44), .B(new_n947), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n952), .ZN(G397));
  OAI211_X1 g528(.A(new_n567), .B(new_n558), .C1(new_n560), .C2(new_n559), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n955));
  AOI22_X1  g530(.A1(new_n571), .A2(KEYINPUT57), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n848), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n482), .A2(new_n490), .B1(new_n957), .B2(new_n487), .ZN(new_n958));
  INV_X1    g533(.A(new_n498), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n497), .B1(new_n482), .B2(new_n494), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n469), .A2(new_n472), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n466), .A2(new_n467), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n965), .B(G40), .C1(new_n966), .C2(new_n463), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n851), .B1(new_n959), .B2(new_n960), .ZN(new_n968));
  INV_X1    g543(.A(new_n850), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n964), .B1(new_n973), .B2(KEYINPUT113), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n971), .B1(new_n852), .B2(new_n962), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(new_n967), .ZN(new_n977));
  AOI21_X1  g552(.A(G1956), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n967), .B1(new_n963), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT106), .B(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT56), .B(G2072), .Z(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n956), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n603), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n967), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n852), .A2(new_n962), .A3(new_n971), .ZN(new_n989));
  AOI21_X1  g564(.A(G1348), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G40), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n468), .A2(new_n473), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n852), .A2(new_n992), .A3(new_n962), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(G2067), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n986), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(KEYINPUT97), .A2(new_n958), .B1(new_n496), .B2(new_n498), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n997), .B2(new_n850), .ZN(new_n998));
  OAI211_X1 g573(.A(KEYINPUT113), .B(new_n992), .C1(new_n998), .C2(new_n971), .ZN(new_n999));
  INV_X1    g574(.A(new_n964), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n977), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1956), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n956), .ZN(new_n1004));
  INV_X1    g579(.A(new_n985), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n996), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n986), .A2(KEYINPUT119), .A3(new_n1006), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT61), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n986), .B2(KEYINPUT119), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n986), .A2(KEYINPUT61), .A3(new_n1006), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n979), .B1(G164), .B2(G1384), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n982), .A2(new_n1013), .A3(new_n1014), .A4(new_n992), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n980), .A2(KEYINPUT117), .A3(new_n1014), .A4(new_n982), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT58), .B(G1341), .Z(new_n1019));
  NAND2_X1  g594(.A1(new_n993), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n547), .B1(new_n1022), .B2(KEYINPUT59), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT118), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1021), .A2(KEYINPUT118), .A3(new_n1025), .A4(new_n548), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n989), .A3(new_n992), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n713), .ZN(new_n1032));
  INV_X1    g607(.A(new_n994), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(KEYINPUT60), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT60), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n990), .A2(new_n1037), .A3(new_n994), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n603), .B1(new_n1038), .B2(KEYINPUT120), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1035), .A3(new_n987), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n995), .A2(KEYINPUT60), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1012), .B(new_n1029), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1007), .B1(new_n1011), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2078), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n980), .A2(new_n1045), .A3(new_n982), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1046), .A2(new_n1047), .B1(new_n1031), .B2(new_n730), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n982), .A2(KEYINPUT53), .A3(new_n1045), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT45), .B1(new_n852), .B2(new_n981), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1050), .A2(KEYINPUT122), .A3(new_n967), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT122), .B1(new_n1050), .B2(new_n967), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(KEYINPUT123), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1055), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1048), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n992), .B1(new_n963), .B2(new_n979), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT45), .B1(new_n852), .B2(new_n962), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(KEYINPUT53), .A3(new_n1045), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1048), .A2(new_n1065), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n1066), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT124), .B1(new_n1066), .B2(G171), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1060), .A2(KEYINPUT54), .A3(new_n1061), .A4(new_n1069), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1064), .A2(G1966), .B1(new_n1031), .B2(G2084), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G286), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1075), .B(G8), .C1(new_n1071), .C2(G286), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(G8), .A3(G286), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n573), .A2(G8), .A3(new_n575), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n573), .A2(KEYINPUT55), .A3(G8), .A4(new_n575), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n999), .A2(new_n977), .A3(new_n708), .A4(new_n1000), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1971), .B1(new_n980), .B2(new_n982), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G8), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT109), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1088), .B(new_n1093), .C1(G2090), .C2(new_n1031), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1031), .A2(G2090), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT109), .B1(new_n1095), .B2(new_n1087), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(new_n1094), .A3(G8), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n507), .A2(G86), .A3(new_n512), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n584), .A2(G651), .B1(G48), .B2(new_n520), .ZN(new_n1101));
  INV_X1    g676(.A(G1981), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT110), .B(new_n1099), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1090), .B1(new_n998), .B2(new_n992), .ZN(new_n1106));
  OAI21_X1  g681(.A(G1981), .B1(new_n581), .B2(new_n587), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(KEYINPUT49), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT110), .B1(new_n1111), .B2(new_n1099), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n578), .B(G1976), .C1(new_n579), .C2(new_n559), .ZN(new_n1114));
  INV_X1    g689(.A(G1976), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(G288), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1106), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n993), .A2(new_n1114), .A3(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT52), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1098), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT110), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(new_n1105), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT114), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1080), .A2(new_n1091), .A3(new_n1097), .A4(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(G301), .B(new_n1048), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1066), .A2(G171), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT54), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1044), .A2(new_n1070), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1125), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NOR4_X1   g710(.A1(new_n1134), .A2(new_n1072), .A3(new_n1135), .A4(G286), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1094), .A2(new_n1096), .A3(G8), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1085), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1097), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1072), .A2(G286), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1127), .A2(new_n1091), .A3(new_n1097), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1108), .B(KEYINPUT111), .ZN(new_n1146));
  NOR2_X1   g721(.A1(G288), .A2(G1976), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT112), .Z(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1148), .B2(new_n1125), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1106), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1097), .A2(new_n1134), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1080), .B(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1127), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n1130), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1133), .A2(new_n1145), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1050), .A2(new_n992), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n723), .A2(new_n1014), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT107), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n761), .B(G2067), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n722), .A2(G1996), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n798), .B(new_n801), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(G290), .B(G1986), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1158), .B1(new_n1162), .B2(new_n863), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT46), .B1(new_n1158), .B2(G1996), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1158), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT47), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n799), .A2(new_n801), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT126), .ZN(new_n1177));
  INV_X1    g752(.A(G2067), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1165), .A2(new_n1177), .B1(new_n1178), .B2(new_n761), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1175), .B1(new_n1179), .B2(new_n1158), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1158), .A2(G1986), .A3(G290), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT48), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1167), .B2(KEYINPUT127), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1167), .A2(KEYINPUT127), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1170), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g761(.A1(G401), .A2(new_n461), .ZN(new_n1188));
  AND4_X1   g762(.A1(new_n662), .A2(new_n684), .A3(new_n685), .A4(new_n1188), .ZN(new_n1189));
  OAI211_X1 g763(.A(new_n875), .B(new_n1189), .C1(new_n941), .C2(new_n944), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


