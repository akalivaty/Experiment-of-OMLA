//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n191));
  OAI211_X1 g005(.A(G119), .B(new_n187), .C1(new_n190), .C2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI22_X1  g007(.A1(new_n188), .A2(new_n189), .B1(new_n193), .B2(G128), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(new_n194), .C1(G119), .C2(new_n187), .ZN(new_n195));
  XNOR2_X1  g009(.A(G119), .B(G128), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT24), .B(G110), .Z(new_n197));
  AOI22_X1  g011(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G140), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT75), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n205), .B2(new_n208), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n198), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n200), .A2(new_n202), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n205), .A2(new_n208), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n213), .B(new_n215), .C1(new_n216), .C2(new_n206), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT22), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G902), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n212), .A2(new_n217), .A3(new_n222), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(G234), .B2(new_n225), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n233));
  INV_X1    g047(.A(new_n231), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n224), .A2(new_n225), .A3(new_n234), .A4(new_n226), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n230), .B1(new_n236), .B2(new_n229), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G143), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n239), .B(G146), .C1(new_n187), .C2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n206), .A2(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n244));
  OAI221_X1 g058(.A(new_n240), .B1(G128), .B2(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G137), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(G137), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n246), .B2(G137), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n252), .A2(new_n254), .A3(new_n255), .A4(new_n247), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n245), .B(new_n250), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT2), .B(G113), .Z(new_n260));
  XNOR2_X1  g074(.A(G116), .B(G119), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  INV_X1    g079(.A(new_n261), .ZN(new_n266));
  INV_X1    g080(.A(new_n260), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n263), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n252), .A2(new_n247), .A3(new_n254), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n241), .A2(new_n242), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G128), .ZN(new_n276));
  XNOR2_X1  g090(.A(G143), .B(G146), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT64), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT64), .B1(new_n243), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n259), .B(new_n268), .C1(new_n273), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n269), .A2(G131), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n257), .B2(new_n258), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n282), .B1(KEYINPUT64), .B2(new_n278), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n268), .B1(new_n293), .B2(new_n259), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n259), .B1(new_n273), .B2(new_n284), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n263), .A2(new_n265), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n267), .A2(new_n266), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(KEYINPUT68), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT28), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n287), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(G101), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n304), .B(new_n306), .Z(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT67), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n285), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n296), .A2(KEYINPUT30), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n259), .B(new_n313), .C1(new_n273), .C2(new_n284), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(new_n299), .ZN(new_n316));
  INV_X1    g130(.A(new_n307), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT31), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n268), .B1(new_n312), .B2(new_n314), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  NOR4_X1   g134(.A1(new_n319), .A2(new_n320), .A3(new_n307), .A4(new_n311), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n310), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G472), .A2(G902), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT32), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n314), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n313), .B1(new_n293), .B2(new_n259), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n299), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n317), .A3(new_n285), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n320), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n328), .A2(KEYINPUT31), .A3(new_n317), .A4(new_n285), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n330), .A2(new_n331), .B1(new_n309), .B2(new_n302), .ZN(new_n332));
  INV_X1    g146(.A(new_n323), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT69), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n322), .A2(new_n335), .A3(new_n323), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n325), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n308), .B(new_n287), .C1(new_n295), .C2(new_n301), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n296), .A2(new_n299), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n288), .A3(new_n285), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT28), .A3(new_n300), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n308), .A4(new_n287), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n307), .B1(new_n319), .B2(new_n311), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n341), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n351), .A3(new_n285), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n296), .A2(KEYINPUT72), .A3(new_n299), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT28), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n287), .A2(KEYINPUT73), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n287), .A2(KEYINPUT73), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n357), .A2(new_n347), .A3(new_n307), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G902), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n340), .B2(KEYINPUT70), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT71), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n346), .A4(new_n348), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n350), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G472), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n238), .B1(new_n339), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(KEYINPUT81), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n292), .A2(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n245), .A2(new_n201), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G224), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G953), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n373), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n377));
  XOR2_X1   g191(.A(G110), .B(G122), .Z(new_n378));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(G104), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n383), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n384));
  OAI22_X1  g198(.A1(new_n383), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n382), .A2(new_n384), .A3(new_n385), .A4(KEYINPUT78), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(G101), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n382), .A2(new_n384), .A3(new_n385), .A4(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n388), .A2(new_n395), .A3(G101), .A4(new_n389), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n299), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n381), .A2(G104), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n383), .A2(G107), .ZN(new_n399));
  OAI21_X1  g213(.A(G101), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n193), .A3(G116), .ZN(new_n404));
  OAI211_X1 g218(.A(G113), .B(new_n404), .C1(new_n266), .C2(new_n403), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n297), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT82), .B1(new_n397), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n378), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n406), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n410), .A2(new_n378), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n377), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n406), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT6), .B1(new_n416), .B2(new_n378), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n376), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n374), .B(new_n375), .C1(KEYINPUT7), .C2(new_n373), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n378), .B(KEYINPUT8), .Z(new_n420));
  INV_X1    g234(.A(new_n406), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n402), .B1(new_n297), .B2(new_n405), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n373), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(new_n411), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n425), .A2(new_n225), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n418), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n418), .B2(new_n426), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n368), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT83), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n418), .A2(new_n426), .ZN(new_n432));
  INV_X1    g246(.A(new_n427), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n418), .A2(new_n426), .A3(new_n427), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n368), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n440));
  INV_X1    g254(.A(G237), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n219), .A3(G214), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n442), .B2(new_n239), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n305), .A2(KEYINPUT86), .A3(G143), .A4(G214), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AND4_X1   g260(.A1(KEYINPUT84), .A2(new_n441), .A3(new_n219), .A4(G214), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT84), .B1(new_n305), .B2(G214), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT85), .B1(new_n449), .B2(new_n239), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n305), .A2(KEYINPUT84), .A3(G214), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n239), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n446), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G131), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT17), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n239), .A3(new_n453), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n454), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n255), .A3(new_n446), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n210), .A2(new_n211), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n255), .B1(new_n462), .B2(new_n446), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n456), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n456), .A2(new_n469), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n215), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(KEYINPUT87), .B(KEYINPUT88), .C1(new_n214), .C2(new_n206), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n214), .A2(new_n206), .ZN(new_n476));
  OR3_X1    g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n470), .A2(new_n471), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n383), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n468), .A2(new_n482), .A3(new_n479), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G475), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n457), .A2(KEYINPUT89), .A3(new_n463), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n492));
  AOI211_X1 g306(.A(G131), .B(new_n445), .C1(new_n461), .C2(new_n454), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n466), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n214), .A2(KEYINPUT90), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT19), .Z(new_n496));
  AOI21_X1  g310(.A(new_n211), .B1(new_n496), .B2(new_n206), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n479), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n490), .B1(new_n499), .B2(new_n483), .ZN(new_n500));
  AOI211_X1 g314(.A(KEYINPUT91), .B(new_n482), .C1(new_n498), .C2(new_n479), .ZN(new_n501));
  INV_X1    g315(.A(new_n485), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G475), .A2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n503), .A2(KEYINPUT20), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n499), .A2(new_n483), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT91), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n499), .A2(new_n490), .A3(new_n483), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n485), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n507), .B1(new_n511), .B2(new_n504), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n489), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G952), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(G953), .ZN(new_n515));
  INV_X1    g329(.A(G234), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(new_n441), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT94), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(G902), .B(G953), .C1(new_n516), .C2(new_n441), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT95), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT21), .B(G898), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n519), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n187), .A2(KEYINPUT92), .A3(G143), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT92), .B1(new_n187), .B2(G143), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT13), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT93), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n187), .A2(G143), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G134), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n246), .A3(new_n530), .ZN(new_n535));
  XNOR2_X1  g349(.A(G116), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n381), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G116), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT14), .A3(G122), .ZN(new_n540));
  INV_X1    g354(.A(new_n536), .ZN(new_n541));
  OAI211_X1 g355(.A(G107), .B(new_n540), .C1(new_n541), .C2(KEYINPUT14), .ZN(new_n542));
  INV_X1    g356(.A(new_n535), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n246), .B1(new_n531), .B2(new_n530), .ZN(new_n544));
  OAI221_X1 g358(.A(new_n542), .B1(G107), .B2(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT9), .B(G234), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n548), .A2(new_n228), .A3(G953), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n538), .A2(new_n545), .A3(new_n549), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n225), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n554), .B(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n513), .A2(new_n525), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G469), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n394), .A2(new_n292), .A3(new_n396), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n402), .A2(KEYINPUT10), .A3(new_n245), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n402), .A2(new_n245), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n560), .A2(new_n273), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n245), .B(new_n401), .Z(new_n566));
  INV_X1    g380(.A(KEYINPUT79), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n291), .ZN(new_n569));
  XNOR2_X1  g383(.A(G110), .B(G140), .ZN(new_n570));
  INV_X1    g384(.A(G227), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G953), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n570), .B(new_n572), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n567), .A2(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n245), .B(new_n401), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n273), .ZN(new_n577));
  AND4_X1   g391(.A1(new_n565), .A2(new_n569), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n291), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n573), .B1(new_n580), .B2(new_n565), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n559), .B(new_n225), .C1(new_n578), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(G469), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n565), .A2(new_n573), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT80), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n565), .A2(new_n586), .A3(new_n573), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n569), .A2(new_n565), .A3(new_n577), .ZN(new_n589));
  INV_X1    g403(.A(new_n573), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n582), .B(new_n583), .C1(new_n592), .C2(new_n559), .ZN(new_n593));
  OAI21_X1  g407(.A(G221), .B1(new_n548), .B2(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n365), .A2(new_n439), .A3(new_n558), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(new_n525), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n368), .B(new_n599), .C1(new_n428), .C2(new_n429), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT20), .B1(new_n503), .B2(new_n505), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n511), .A2(new_n507), .A3(new_n504), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n488), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n550), .B2(KEYINPUT96), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n553), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n551), .A2(new_n552), .A3(new_n605), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n555), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n554), .A2(G478), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n555), .A2(new_n225), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n600), .A2(new_n603), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n596), .A2(new_n237), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n322), .B2(new_n225), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n337), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND3_X1  g437(.A1(new_n601), .A2(KEYINPUT97), .A3(new_n602), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n486), .B2(new_n487), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n482), .B1(new_n468), .B2(new_n479), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n225), .B1(new_n502), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT98), .A3(G475), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n511), .A2(new_n631), .A3(new_n507), .A4(new_n504), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n624), .A2(new_n557), .A3(new_n630), .A4(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n600), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n620), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G107), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT99), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(G9));
  NAND2_X1  g453(.A1(new_n236), .A2(new_n229), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n218), .B(KEYINPUT100), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n223), .A2(KEYINPUT36), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n641), .B(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n225), .B1(new_n228), .B2(G234), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n337), .A2(new_n618), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n439), .A2(new_n558), .A3(new_n596), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT37), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(G110), .Z(G12));
  INV_X1    g465(.A(new_n646), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n339), .B2(new_n364), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n519), .B1(new_n654), .B2(new_n522), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n593), .A2(new_n594), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n430), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n653), .A2(new_n634), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  NAND2_X1  g474(.A1(new_n352), .A2(new_n353), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n329), .B1(new_n308), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n225), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n339), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n655), .B(KEYINPUT39), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n595), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n339), .A2(new_n670), .A3(new_n664), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n513), .A2(new_n652), .A3(new_n368), .A4(new_n557), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n436), .B(KEYINPUT38), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n672), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n239), .ZN(G45));
  NOR3_X1   g494(.A1(new_n603), .A2(new_n613), .A3(new_n657), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n337), .A2(new_n338), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n364), .A2(new_n682), .A3(new_n324), .ZN(new_n683));
  INV_X1    g497(.A(new_n430), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n683), .A3(new_n684), .A4(new_n646), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NOR2_X1   g500(.A1(new_n578), .A2(new_n581), .ZN(new_n687));
  OAI21_X1  g501(.A(G469), .B1(new_n687), .B2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n582), .ZN(new_n689));
  INV_X1    g503(.A(new_n594), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n365), .A2(new_n614), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n365), .A2(new_n634), .A3(new_n635), .A4(new_n691), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT103), .B(G116), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G18));
  OAI211_X1 g511(.A(new_n691), .B(new_n368), .C1(new_n428), .C2(new_n429), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n653), .A2(new_n558), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  INV_X1    g515(.A(new_n557), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n603), .A2(new_n430), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n330), .A2(new_n331), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n357), .A2(new_n309), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n333), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n617), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n238), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n703), .A2(new_n599), .A3(new_n691), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NOR3_X1   g525(.A1(new_n603), .A2(new_n613), .A3(new_n655), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n652), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n699), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  NAND3_X1  g529(.A1(new_n434), .A2(new_n368), .A3(new_n435), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n322), .A2(new_n323), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT104), .B1(new_n719), .B2(new_n338), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n333), .B1(new_n704), .B2(new_n310), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(KEYINPUT32), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n332), .A2(KEYINPUT105), .A3(new_n338), .A4(new_n333), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n722), .B2(KEYINPUT32), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n324), .A2(KEYINPUT105), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n722), .A2(new_n721), .A3(KEYINPUT32), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n725), .A2(new_n730), .A3(new_n364), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n237), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n731), .B2(new_n237), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n681), .B(new_n718), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n615), .B1(new_n339), .B2(new_n364), .ZN(new_n736));
  INV_X1    g550(.A(new_n716), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n712), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n717), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND4_X1  g556(.A1(new_n736), .A2(new_n634), .A3(new_n656), .A4(new_n737), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT107), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n246), .ZN(G36));
  OAI211_X1 g559(.A(new_n612), .B(new_n489), .C1(new_n506), .C2(new_n512), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT43), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n603), .A2(new_n748), .A3(new_n612), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n749), .A3(new_n619), .A4(new_n646), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n592), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n588), .A2(KEYINPUT45), .A3(new_n591), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n583), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n583), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n582), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n594), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n667), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n716), .B(KEYINPUT108), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n750), .B2(new_n751), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n253), .ZN(G39));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n594), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n683), .A2(new_n237), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n712), .A3(new_n737), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NOR2_X1   g589(.A1(new_n733), .A2(new_n734), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n747), .A2(new_n519), .A3(new_n749), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n691), .A2(new_n434), .A3(new_n368), .A4(new_n435), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT48), .Z(new_n783));
  AND2_X1   g597(.A1(new_n666), .A2(new_n671), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n518), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n603), .A2(new_n613), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n237), .A3(new_n786), .A4(new_n780), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n747), .A2(new_n709), .A3(new_n749), .A4(new_n519), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n699), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n783), .A2(new_n515), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n691), .A2(new_n367), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n788), .A2(new_n676), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT50), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n513), .A2(new_n612), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n785), .A2(new_n237), .A3(new_n797), .A4(new_n780), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n777), .A2(new_n713), .A3(new_n780), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT117), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n789), .A2(KEYINPUT114), .A3(new_n765), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT114), .B1(new_n789), .B2(new_n765), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n689), .A2(new_n594), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n801), .A2(new_n802), .B1(new_n772), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n796), .A2(new_n798), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n806), .A3(KEYINPUT51), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n791), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n698), .A2(new_n603), .A3(new_n613), .A4(new_n655), .ZN(new_n812));
  INV_X1    g626(.A(new_n657), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n436), .A2(new_n813), .A3(new_n368), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n633), .A2(new_n814), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n812), .A2(new_n713), .B1(new_n815), .B2(new_n653), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n603), .A2(new_n702), .A3(new_n646), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n665), .A3(new_n658), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(KEYINPUT52), .A3(new_n685), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n659), .A2(new_n685), .A3(new_n714), .A4(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(KEYINPUT112), .A3(new_n821), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n695), .A2(new_n692), .A3(new_n710), .A4(new_n700), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n557), .B(new_n489), .C1(new_n506), .C2(new_n512), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n603), .B2(new_n613), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n439), .A2(new_n829), .A3(new_n599), .A4(new_n620), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n597), .A2(new_n649), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n708), .A2(new_n603), .A3(new_n613), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n624), .A2(new_n630), .A3(new_n632), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n339), .B2(new_n364), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n835), .B2(new_n702), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n737), .A2(new_n646), .A3(new_n813), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT110), .B(new_n743), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n839));
  INV_X1    g653(.A(new_n743), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n630), .A2(new_n632), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n506), .A2(new_n512), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(KEYINPUT97), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n683), .A2(new_n843), .A3(new_n702), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n786), .A2(new_n707), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n837), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n832), .A2(new_n741), .A3(new_n838), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n847), .A2(new_n838), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n819), .A2(new_n822), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n741), .A3(new_n852), .A4(new_n832), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n826), .A2(new_n850), .B1(new_n853), .B2(new_n849), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n853), .A2(new_n849), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n851), .A2(new_n858), .A3(new_n741), .A4(new_n832), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n848), .A2(KEYINPUT111), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n826), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n857), .B1(new_n861), .B2(new_n849), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n811), .B(new_n856), .C1(new_n855), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n514), .A2(new_n219), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n746), .A2(new_n367), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n238), .B1(new_n689), .B2(KEYINPUT49), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n594), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT109), .Z(new_n869));
  NOR2_X1   g683(.A1(new_n689), .A2(KEYINPUT49), .ZN(new_n870));
  OR4_X1    g684(.A1(new_n676), .A2(new_n869), .A3(new_n784), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n871), .ZN(G75));
  NAND2_X1  g686(.A1(new_n514), .A2(G953), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n826), .ZN(new_n875));
  INV_X1    g689(.A(new_n852), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n849), .B1(new_n848), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n225), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n412), .A2(new_n417), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n376), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n874), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT118), .B1(new_n854), .B2(new_n225), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n875), .A2(new_n877), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(G902), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n888), .A3(new_n433), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n884), .B1(new_n889), .B2(new_n891), .ZN(G51));
  INV_X1    g706(.A(new_n874), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n583), .B(KEYINPUT57), .Z(new_n894));
  AND3_X1   g708(.A1(new_n875), .A2(new_n855), .A3(new_n877), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n855), .B1(new_n875), .B2(new_n877), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n687), .B(KEYINPUT121), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n756), .B(KEYINPUT122), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n885), .A2(new_n888), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n899), .B2(new_n901), .ZN(G54));
  AND2_X1   g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n885), .A2(new_n888), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n511), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n885), .A2(new_n888), .A3(new_n503), .A4(new_n903), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n893), .B1(new_n905), .B2(new_n906), .ZN(G60));
  AND2_X1   g721(.A1(new_n607), .A2(new_n608), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n856), .B1(new_n862), .B2(new_n855), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n611), .B(KEYINPUT59), .Z(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n908), .B(new_n910), .C1(new_n895), .C2(new_n896), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n874), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(G63));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n854), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n224), .A2(new_n226), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n874), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n917), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n886), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n644), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n915), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n893), .B1(new_n923), .B2(new_n919), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n926), .B(KEYINPUT61), .C1(new_n644), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(G66));
  OAI21_X1  g742(.A(G953), .B1(new_n524), .B2(new_n372), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n832), .B2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n880), .B1(G898), .B2(new_n219), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(G69));
  OAI21_X1  g746(.A(G953), .B1(new_n571), .B2(new_n654), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n763), .B(new_n703), .C1(new_n733), .C2(new_n734), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n741), .A2(new_n774), .A3(new_n743), .A4(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n659), .A2(new_n685), .A3(new_n714), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n764), .B2(new_n766), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n937), .B(KEYINPUT124), .C1(new_n764), .C2(new_n766), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(G953), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n315), .B(new_n496), .Z(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n816), .A2(new_n685), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n679), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n675), .A2(new_n676), .ZN(new_n949));
  INV_X1    g763(.A(new_n678), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n784), .A3(new_n950), .A4(new_n669), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(KEYINPUT62), .A3(new_n937), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n774), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n767), .ZN(new_n955));
  INV_X1    g769(.A(new_n829), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n738), .A2(new_n667), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n959), .A2(new_n219), .A3(new_n944), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n934), .B1(new_n945), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n654), .B1(new_n944), .B2(new_n571), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n219), .B2(new_n962), .ZN(G72));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n316), .B(KEYINPUT125), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n307), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n940), .A2(new_n941), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n741), .A2(new_n774), .A3(new_n743), .A4(new_n935), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n832), .ZN(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT126), .B1(new_n972), .B2(new_n893), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n974));
  INV_X1    g788(.A(new_n971), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n942), .B2(new_n832), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n974), .B(new_n874), .C1(new_n976), .C2(new_n966), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n953), .A2(new_n955), .A3(new_n832), .A4(new_n958), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n965), .B1(new_n979), .B2(new_n971), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n317), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n975), .B1(new_n348), .B2(new_n329), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n862), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n964), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n307), .B(new_n965), .C1(new_n979), .C2(new_n971), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n861), .A2(new_n849), .ZN(new_n987));
  INV_X1    g801(.A(new_n857), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n986), .B1(new_n989), .B2(new_n982), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(KEYINPUT127), .A3(new_n973), .A4(new_n977), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n985), .A2(new_n991), .ZN(G57));
endmodule


