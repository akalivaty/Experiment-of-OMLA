

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  NOR2_X2 U323 ( .A1(n463), .A2(n529), .ZN(n571) );
  NOR2_X1 U324 ( .A1(n557), .A2(n576), .ZN(n369) );
  XNOR2_X1 U325 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U326 ( .A(n435), .B(n337), .ZN(n340) );
  INV_X1 U327 ( .A(KEYINPUT48), .ZN(n400) );
  XNOR2_X1 U328 ( .A(n401), .B(n400), .ZN(n551) );
  XOR2_X1 U329 ( .A(n348), .B(n347), .Z(n581) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n465) );
  XNOR2_X1 U331 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U332 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n447) );
  XOR2_X1 U334 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n292) );
  NAND2_X1 U335 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n299) );
  INV_X1 U337 ( .A(G218GAT), .ZN(n293) );
  NAND2_X1 U338 ( .A1(KEYINPUT80), .A2(n293), .ZN(n296) );
  INV_X1 U339 ( .A(KEYINPUT80), .ZN(n294) );
  NAND2_X1 U340 ( .A1(n294), .A2(G218GAT), .ZN(n295) );
  NAND2_X1 U341 ( .A1(n296), .A2(n295), .ZN(n298) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n372) );
  XOR2_X1 U344 ( .A(n299), .B(n372), .Z(n302) );
  XNOR2_X1 U345 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n300), .B(G211GAT), .ZN(n434) );
  XNOR2_X1 U347 ( .A(G8GAT), .B(n434), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(G176GAT), .B(G64GAT), .Z(n344) );
  XOR2_X1 U350 ( .A(n303), .B(n344), .Z(n305) );
  XNOR2_X1 U351 ( .A(G204GAT), .B(G92GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U353 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n307) );
  XNOR2_X1 U354 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(G169GAT), .B(n308), .Z(n462) );
  XNOR2_X1 U357 ( .A(n309), .B(n462), .ZN(n470) );
  INV_X1 U358 ( .A(n470), .ZN(n526) );
  XOR2_X1 U359 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n392) );
  XOR2_X1 U360 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n311) );
  XNOR2_X1 U361 ( .A(G127GAT), .B(G64GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n326) );
  XOR2_X1 U363 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XOR2_X1 U364 ( .A(G211GAT), .B(G78GAT), .Z(n313) );
  XNOR2_X1 U365 ( .A(G183GAT), .B(G71GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n440), .B(n314), .Z(n316) );
  NAND2_X1 U368 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U370 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n324) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G8GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n321), .B(G1GAT), .ZN(n361) );
  XNOR2_X1 U376 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n322), .B(KEYINPUT74), .ZN(n339) );
  XNOR2_X1 U378 ( .A(n361), .B(n339), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n572) );
  XOR2_X1 U381 ( .A(KEYINPUT77), .B(G92GAT), .Z(n328) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G85GAT), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U384 ( .A(G106GAT), .B(n329), .Z(n379) );
  XOR2_X1 U385 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n331) );
  XNOR2_X1 U386 ( .A(KEYINPUT75), .B(KEYINPUT78), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n379), .B(n332), .ZN(n348) );
  XOR2_X1 U389 ( .A(G78GAT), .B(G148GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(KEYINPUT76), .B(G204GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n435) );
  NAND2_X1 U392 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  INV_X1 U393 ( .A(KEYINPUT33), .ZN(n335) );
  INV_X1 U394 ( .A(n340), .ZN(n338) );
  NAND2_X1 U395 ( .A1(n338), .A2(n339), .ZN(n343) );
  INV_X1 U396 ( .A(n339), .ZN(n341) );
  NAND2_X1 U397 ( .A1(n341), .A2(n340), .ZN(n342) );
  NAND2_X1 U398 ( .A1(n343), .A2(n342), .ZN(n346) );
  XOR2_X1 U399 ( .A(G120GAT), .B(G71GAT), .Z(n451) );
  XNOR2_X1 U400 ( .A(n451), .B(n344), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U402 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n581), .B(n349), .ZN(n566) );
  INV_X1 U404 ( .A(n566), .ZN(n557) );
  XOR2_X1 U405 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n351) );
  XNOR2_X1 U406 ( .A(KEYINPUT70), .B(KEYINPUT73), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n368) );
  XOR2_X1 U408 ( .A(G197GAT), .B(G22GAT), .Z(n353) );
  XNOR2_X1 U409 ( .A(G36GAT), .B(G50GAT), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U411 ( .A(KEYINPUT30), .B(G113GAT), .Z(n355) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G141GAT), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U414 ( .A(n357), .B(n356), .Z(n366) );
  XOR2_X1 U415 ( .A(KEYINPUT7), .B(KEYINPUT72), .Z(n359) );
  XNOR2_X1 U416 ( .A(G43GAT), .B(G29GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U418 ( .A(KEYINPUT8), .B(n360), .Z(n389) );
  XOR2_X1 U419 ( .A(n361), .B(KEYINPUT71), .Z(n363) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n389), .B(n364), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(n368), .B(n367), .Z(n564) );
  INV_X1 U425 ( .A(n564), .ZN(n576) );
  XNOR2_X1 U426 ( .A(n369), .B(KEYINPUT46), .ZN(n370) );
  NOR2_X1 U427 ( .A1(n572), .A2(n370), .ZN(n390) );
  XOR2_X1 U428 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  INV_X1 U429 ( .A(n441), .ZN(n371) );
  NAND2_X1 U430 ( .A1(n372), .A2(n371), .ZN(n375) );
  INV_X1 U431 ( .A(n372), .ZN(n373) );
  NAND2_X1 U432 ( .A1(n373), .A2(n441), .ZN(n374) );
  NAND2_X1 U433 ( .A1(n375), .A2(n374), .ZN(n377) );
  NAND2_X1 U434 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U437 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n381) );
  XNOR2_X1 U438 ( .A(G134GAT), .B(KEYINPUT79), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U440 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n383) );
  XNOR2_X1 U441 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U443 ( .A(n385), .B(n384), .Z(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n393) );
  NAND2_X1 U446 ( .A1(n390), .A2(n393), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n399) );
  XNOR2_X1 U448 ( .A(KEYINPUT81), .B(n393), .ZN(n464) );
  INV_X1 U449 ( .A(n464), .ZN(n547) );
  XNOR2_X1 U450 ( .A(n547), .B(KEYINPUT36), .ZN(n590) );
  INV_X1 U451 ( .A(n572), .ZN(n585) );
  NOR2_X1 U452 ( .A1(n590), .A2(n585), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n394), .B(KEYINPUT45), .ZN(n395) );
  NAND2_X1 U454 ( .A1(n395), .A2(n581), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n396), .B(KEYINPUT115), .ZN(n397) );
  NAND2_X1 U456 ( .A1(n397), .A2(n576), .ZN(n398) );
  NAND2_X1 U457 ( .A1(n399), .A2(n398), .ZN(n401) );
  NOR2_X1 U458 ( .A1(n526), .A2(n551), .ZN(n402) );
  XNOR2_X1 U459 ( .A(KEYINPUT54), .B(n402), .ZN(n427) );
  XOR2_X1 U460 ( .A(G57GAT), .B(G148GAT), .Z(n404) );
  XNOR2_X1 U461 ( .A(G1GAT), .B(G120GAT), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G155GAT), .Z(n406) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G162GAT), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n426) );
  XOR2_X1 U467 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT4), .B(KEYINPUT97), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U470 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n412) );
  XNOR2_X1 U471 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U473 ( .A(n414), .B(n413), .Z(n424) );
  XNOR2_X1 U474 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n415), .B(KEYINPUT87), .ZN(n416) );
  XOR2_X1 U476 ( .A(n416), .B(KEYINPUT86), .Z(n418) );
  XNOR2_X1 U477 ( .A(G113GAT), .B(G134GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n458) );
  XNOR2_X1 U479 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n419), .B(KEYINPUT2), .ZN(n438) );
  XOR2_X1 U481 ( .A(KEYINPUT96), .B(n438), .Z(n421) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n458), .B(n422), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n523) );
  NAND2_X1 U487 ( .A1(n427), .A2(n523), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n428), .B(KEYINPUT65), .ZN(n575) );
  XOR2_X1 U489 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n430) );
  XNOR2_X1 U490 ( .A(G218GAT), .B(G106GAT), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n445) );
  XOR2_X1 U492 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n432) );
  NAND2_X1 U493 ( .A1(G228GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U495 ( .A(n433), .B(KEYINPUT23), .Z(n437) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n474) );
  NAND2_X1 U502 ( .A1(n575), .A2(n474), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n463) );
  XOR2_X1 U504 ( .A(KEYINPUT89), .B(G176GAT), .Z(n449) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(G99GAT), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U507 ( .A(n450), .B(G190GAT), .Z(n453) );
  XNOR2_X1 U508 ( .A(G43GAT), .B(n451), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n455) );
  NAND2_X1 U511 ( .A1(G227GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U513 ( .A(n457), .B(n456), .Z(n460) );
  XNOR2_X1 U514 ( .A(n458), .B(KEYINPUT88), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n529) );
  NAND2_X1 U517 ( .A1(n571), .A2(n464), .ZN(n468) );
  XOR2_X1 U518 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n466) );
  AND2_X1 U519 ( .A1(n581), .A2(n564), .ZN(n498) );
  INV_X1 U520 ( .A(n529), .ZN(n538) );
  XOR2_X1 U521 ( .A(n526), .B(KEYINPUT27), .Z(n477) );
  INV_X1 U522 ( .A(n523), .ZN(n553) );
  XNOR2_X1 U523 ( .A(n474), .B(KEYINPUT28), .ZN(n532) );
  AND2_X1 U524 ( .A1(n553), .A2(n532), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n477), .A2(n469), .ZN(n536) );
  NOR2_X1 U526 ( .A1(n538), .A2(n536), .ZN(n482) );
  NAND2_X1 U527 ( .A1(n470), .A2(n538), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n471), .A2(n474), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT25), .ZN(n478) );
  XNOR2_X1 U531 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n538), .A2(n474), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(n574) );
  NAND2_X1 U534 ( .A1(n574), .A2(n477), .ZN(n550) );
  NAND2_X1 U535 ( .A1(n478), .A2(n550), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n523), .A2(n479), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT102), .B(n480), .Z(n481) );
  NOR2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n495) );
  XOR2_X1 U539 ( .A(KEYINPUT85), .B(KEYINPUT16), .Z(n484) );
  NAND2_X1 U540 ( .A1(n572), .A2(n547), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n495), .A2(n485), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT103), .B(n486), .Z(n510) );
  NAND2_X1 U544 ( .A1(n498), .A2(n510), .ZN(n493) );
  NOR2_X1 U545 ( .A1(n523), .A2(n493), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U548 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  NOR2_X1 U549 ( .A1(n526), .A2(n493), .ZN(n490) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n490), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n529), .A2(n493), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n532), .A2(n493), .ZN(n494) );
  XOR2_X1 U555 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  NOR2_X1 U556 ( .A1(n590), .A2(n495), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n585), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n497), .ZN(n522) );
  NAND2_X1 U559 ( .A1(n498), .A2(n522), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT38), .ZN(n507) );
  NOR2_X1 U561 ( .A1(n523), .A2(n507), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n500), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT39), .ZN(G1328GAT) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n503) );
  NOR2_X1 U565 ( .A1(n526), .A2(n507), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n507), .A2(n529), .ZN(n505) );
  XNOR2_X1 U568 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U570 ( .A(G43GAT), .B(n506), .Z(G1330GAT) );
  NOR2_X1 U571 ( .A1(n507), .A2(n532), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  NOR2_X1 U574 ( .A1(n564), .A2(n557), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n510), .A2(n521), .ZN(n517) );
  NOR2_X1 U576 ( .A1(n523), .A2(n517), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n517), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n529), .A2(n517), .ZN(n516) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n532), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n531) );
  NOR2_X1 U590 ( .A1(n523), .A2(n531), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n531), .ZN(n527) );
  XOR2_X1 U594 ( .A(KEYINPUT112), .B(n527), .Z(n528) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n531), .ZN(n530) );
  XOR2_X1 U597 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U599 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n551), .A2(n536), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n546) );
  NOR2_X1 U604 ( .A1(n576), .A2(n546), .ZN(n539) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n557), .A2(n546), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n585), .A2(n546), .ZN(n544) );
  XNOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT118), .ZN(n562) );
  NOR2_X1 U620 ( .A1(n562), .A2(n576), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XNOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n557), .A2(n562), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n585), .A2(n562), .ZN(n561) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n393), .ZN(n563) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n571), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT121), .Z(n568) );
  NAND2_X1 U634 ( .A1(n571), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n589) );
  NOR2_X1 U641 ( .A1(n589), .A2(n576), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n589), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n589), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT125), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

