//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n221), .B1(new_n203), .B2(new_n222), .C1(new_n206), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n212), .B1(new_n216), .B2(new_n220), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n213), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n202), .A2(new_n214), .ZN(new_n250));
  XOR2_X1   g0050(.A(KEYINPUT8), .B(G58), .Z(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n214), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n249), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n249), .B1(new_n259), .B2(G20), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G50), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT71), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT67), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G222), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(new_n203), .C2(new_n277), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI211_X1 g0087(.A(G1), .B(G13), .C1(new_n273), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(new_n290), .B2(G226), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n266), .A2(new_n267), .B1(G190), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n265), .A2(KEYINPUT9), .B1(G200), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n294), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT67), .B1(new_n268), .B2(new_n269), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n274), .A2(new_n271), .A3(new_n275), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G107), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n302), .A2(new_n303), .A3(G232), .A4(new_n278), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(G238), .A4(G1698), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT68), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT68), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n305), .A2(new_n310), .A3(new_n306), .A4(new_n307), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n282), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT69), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n286), .B1(new_n290), .B2(G244), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n301), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT69), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n253), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n251), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(KEYINPUT70), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(KEYINPUT70), .B2(new_n325), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n249), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n260), .A2(G77), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n262), .B2(G77), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n317), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n264), .B1(new_n293), .B2(G169), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n301), .B2(new_n293), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n300), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n262), .A2(G68), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT12), .ZN(new_n338));
  INV_X1    g0138(.A(new_n260), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n218), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n218), .A2(G20), .ZN(new_n343));
  INV_X1    g0143(.A(G50), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n343), .B1(new_n253), .B2(new_n203), .C1(new_n256), .C2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n345), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT11), .B1(new_n345), .B2(new_n249), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n286), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n288), .A2(G238), .A3(new_n284), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT73), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT73), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n302), .A2(new_n303), .A3(G232), .A4(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n277), .A2(new_n359), .A3(G226), .A4(new_n278), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n302), .A2(new_n303), .A3(G226), .A4(new_n278), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT72), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n355), .B1(new_n363), .B2(new_n288), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(new_n358), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n361), .A2(KEYINPUT72), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n361), .A2(KEYINPUT72), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n282), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n355), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n372), .A3(G179), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT74), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n373), .B(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n371), .B1(new_n370), .B2(new_n355), .ZN(new_n376));
  AOI211_X1 g0176(.A(KEYINPUT13), .B(new_n354), .C1(new_n369), .C2(new_n282), .ZN(new_n377));
  OAI21_X1  g0177(.A(G169), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n365), .A2(new_n372), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(G169), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n349), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n348), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n365), .B2(new_n372), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n214), .B1(new_n219), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(KEYINPUT76), .B1(G159), .B2(new_n255), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n219), .A2(new_n391), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G20), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n275), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT75), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n268), .B2(new_n269), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n274), .A2(KEYINPUT75), .A3(new_n275), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n214), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n398), .B(KEYINPUT16), .C1(new_n406), .C2(new_n218), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n393), .A2(new_n397), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n302), .B2(new_n303), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n399), .B1(new_n409), .B2(KEYINPUT7), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n410), .B2(G68), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n407), .B(new_n249), .C1(new_n411), .C2(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n252), .B1(new_n259), .B2(G20), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n339), .A2(new_n249), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n413), .A2(new_n414), .B1(new_n339), .B2(new_n252), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n274), .A2(new_n275), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n278), .A2(G226), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(G223), .C2(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n288), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G232), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n350), .B1(new_n289), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G169), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(G179), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n412), .A2(new_n415), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT18), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n420), .A2(new_n386), .A3(new_n422), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n424), .B2(G200), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n412), .A2(new_n415), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT17), .ZN(new_n432));
  OAI21_X1  g0232(.A(G190), .B1(new_n315), .B2(new_n316), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n319), .A2(G200), .A3(new_n321), .ZN(new_n434));
  INV_X1    g0234(.A(new_n331), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n336), .A2(new_n385), .A3(new_n390), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n339), .A2(new_n206), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT25), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT84), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n339), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT83), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n248), .A2(new_n213), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(new_n260), .C1(G1), .C2(new_n273), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n442), .A2(new_n444), .B1(G107), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT23), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n214), .B2(G107), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G87), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n455), .A2(KEYINPUT22), .A3(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n302), .A2(new_n303), .A3(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n214), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT22), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT24), .B(new_n454), .C1(new_n459), .C2(new_n457), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n249), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n448), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n470), .A2(new_n282), .A3(new_n285), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n470), .A2(G264), .A3(new_n288), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G294), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n273), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G250), .A2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(G1698), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(new_n416), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n282), .B1(new_n480), .B2(KEYINPUT85), .ZN(new_n481));
  INV_X1    g0281(.A(G250), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n278), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(G1698), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n484), .C1(new_n268), .C2(new_n269), .ZN(new_n485));
  INV_X1    g0285(.A(new_n476), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT85), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n472), .B(new_n474), .C1(new_n481), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G169), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT86), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n493), .A3(G169), .ZN(new_n494));
  INV_X1    g0294(.A(new_n490), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G179), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n490), .A2(new_n498), .A3(new_n388), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n499), .A2(new_n464), .A3(new_n448), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n498), .B1(new_n490), .B2(new_n388), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G190), .B2(new_n490), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n465), .A2(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n260), .A2(G97), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n447), .B2(G97), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n508), .A2(new_n205), .A3(G107), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n214), .B1(new_n270), .B2(new_n276), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n400), .B1(new_n514), .B2(new_n405), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n515), .B2(new_n206), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n506), .B1(new_n516), .B2(new_n249), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(new_n278), .C1(new_n268), .C2(new_n269), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n518), .A2(new_n519), .B1(G33), .B2(G283), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n302), .A2(new_n303), .A3(G250), .A4(G1698), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n519), .A2(new_n222), .A3(G1698), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n302), .A2(new_n303), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n282), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n470), .A2(G257), .A3(new_n288), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n470), .A2(KEYINPUT77), .A3(G257), .A4(new_n288), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n471), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(G190), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n530), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n517), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n255), .A2(G77), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n510), .B1(new_n508), .B2(new_n507), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(new_n214), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n410), .B2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n505), .B1(new_n538), .B2(new_n445), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n525), .A2(G179), .A3(new_n530), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n320), .B1(new_n525), .B2(new_n530), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n467), .A2(new_n482), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n288), .B1(G274), .B2(new_n467), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G238), .A2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n222), .B2(G1698), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n416), .B1(G33), .B2(G116), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n288), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  OAI211_X1 g0353(.A(G190), .B(new_n548), .C1(new_n551), .C2(new_n288), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n214), .B1(new_n357), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G87), .B2(new_n207), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n214), .B(G68), .C1(new_n268), .C2(new_n269), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n555), .B1(new_n253), .B2(new_n205), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n249), .B1(new_n339), .B2(new_n323), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n447), .A2(G87), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n553), .A2(new_n554), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n249), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n323), .A2(new_n339), .ZN(new_n565));
  INV_X1    g0365(.A(new_n323), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n414), .B(new_n566), .C1(G1), .C2(new_n273), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n552), .A2(new_n320), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n301), .B(new_n548), .C1(new_n551), .C2(new_n288), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n563), .A2(new_n571), .A3(KEYINPUT79), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n503), .A2(new_n544), .A3(new_n546), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n223), .A2(G1698), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n416), .B(new_n578), .C1(G257), .C2(G1698), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G303), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n302), .B2(new_n303), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n282), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n470), .A2(new_n288), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n471), .B1(G270), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G169), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT81), .ZN(new_n589));
  AOI21_X1  g0389(.A(G20), .B1(new_n273), .B2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(G283), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n273), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G116), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G20), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n249), .A2(KEYINPUT80), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT80), .B1(new_n249), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT20), .B(new_n592), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n339), .A2(new_n593), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n446), .B2(new_n593), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n589), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT81), .B(new_n603), .C1(new_n599), .C2(new_n600), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n588), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n601), .A2(new_n604), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n601), .A2(new_n589), .A3(new_n604), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n586), .A2(new_n301), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n588), .B(KEYINPUT21), .C1(new_n605), .C2(new_n606), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n586), .A2(G200), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n585), .A2(new_n583), .A3(G190), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n611), .A2(new_n612), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n609), .A2(new_n615), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n587), .B1(new_n611), .B2(new_n612), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n623), .A2(KEYINPUT21), .B1(new_n613), .B2(new_n614), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT82), .A3(new_n609), .A4(new_n619), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n577), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n438), .A2(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n432), .ZN(new_n628));
  INV_X1    g0428(.A(new_n390), .ZN(new_n629));
  INV_X1    g0429(.A(new_n332), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(new_n384), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  INV_X1    g0433(.A(new_n428), .ZN(new_n634));
  OR3_X1    g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n300), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n335), .ZN(new_n638));
  INV_X1    g0438(.A(new_n571), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n532), .A2(G169), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n301), .B2(new_n532), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n574), .A2(new_n641), .A3(new_n539), .A4(new_n575), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT89), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n517), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n561), .A2(new_n562), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n550), .A2(new_n416), .ZN(new_n648));
  NAND2_X1  g0448(.A1(G33), .A2(G116), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n288), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n548), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n647), .B1(G190), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n552), .A2(new_n654), .A3(G200), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n552), .B2(G200), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n639), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n640), .B(KEYINPUT89), .C1(new_n301), .C2(new_n532), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n645), .A2(new_n646), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n546), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n545), .B1(new_n534), .B2(new_n542), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n659), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n502), .B2(new_n500), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n497), .A2(new_n465), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(new_n609), .A3(new_n616), .A4(new_n615), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n438), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n638), .A2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n259), .A2(new_n214), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT91), .Z(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G343), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n611), .B2(new_n612), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n622), .B2(new_n625), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n624), .A2(new_n609), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n679), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n465), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n503), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n668), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n687), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n682), .A2(new_n679), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n695), .A2(new_n503), .B1(new_n690), .B2(new_n679), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  NOR3_X1   g0497(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT92), .Z(new_n699));
  INV_X1    g0499(.A(new_n210), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n699), .A2(new_n259), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n220), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  AND2_X1   g0505(.A1(new_n525), .A2(new_n530), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n495), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n652), .A2(G179), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(KEYINPUT94), .A3(new_n586), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT94), .B1(new_n708), .B2(new_n586), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n474), .B1(new_n481), .B2(new_n489), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n552), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n614), .A2(new_n713), .A3(new_n706), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n716), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n614), .A2(new_n713), .A3(new_n706), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n711), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n687), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n626), .B2(new_n679), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT95), .B1(new_n726), .B2(new_n685), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n622), .A2(new_n625), .ZN(new_n728));
  INV_X1    g0528(.A(new_n577), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n679), .ZN(new_n730));
  INV_X1    g0530(.A(new_n725), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT95), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n687), .B1(new_n662), .B2(new_n670), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n644), .B1(new_n540), .B2(new_n541), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n659), .A2(new_n660), .A3(new_n539), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT26), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n571), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n740), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT97), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n544), .A2(new_n747), .A3(new_n546), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT97), .B1(new_n663), .B2(new_n664), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n669), .A4(new_n667), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(new_n743), .A3(KEYINPUT96), .A4(new_n571), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n739), .B1(new_n753), .B2(new_n679), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n738), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n735), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n705), .B1(new_n757), .B2(G1), .ZN(G364));
  OAI211_X1 g0558(.A(G1), .B(G13), .C1(new_n214), .C2(G169), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(KEYINPUT99), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n386), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n214), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G294), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n301), .A2(new_n388), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n214), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(KEYINPUT33), .A2(G317), .ZN(new_n771));
  AND2_X1   g0571(.A1(KEYINPUT33), .A2(G317), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n768), .A2(new_n301), .A3(new_n388), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G329), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n766), .A2(new_n773), .A3(new_n304), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n301), .A2(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(new_n768), .A3(KEYINPUT100), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(KEYINPUT100), .B1(new_n778), .B2(new_n768), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n214), .A2(new_n386), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n778), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n388), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n768), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n786), .A2(new_n787), .B1(new_n789), .B2(new_n591), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(new_n767), .ZN(new_n791));
  INV_X1    g0591(.A(G326), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n785), .A2(new_n788), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n581), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n777), .A2(new_n784), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT101), .ZN(new_n796));
  INV_X1    g0596(.A(new_n791), .ZN(new_n797));
  INV_X1    g0597(.A(new_n786), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G50), .A2(new_n797), .B1(new_n798), .B2(G58), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n765), .A2(G97), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n799), .A2(new_n277), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n789), .A2(new_n206), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n793), .A2(new_n455), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(G68), .C2(new_n770), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n774), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n782), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n801), .B(new_n808), .C1(G77), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n762), .B1(new_n796), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n762), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n402), .A2(new_n403), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n700), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G45), .B2(new_n220), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G45), .B2(new_n246), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n304), .A2(new_n700), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(G355), .B(KEYINPUT98), .Z(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n822), .B1(G116), .B2(new_n210), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n815), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n214), .A2(G13), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n259), .B1(new_n825), .B2(G45), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n701), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n811), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n684), .B2(new_n814), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n686), .A2(new_n828), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n684), .A2(new_n685), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  AND4_X1   g0634(.A1(new_n322), .A2(new_n317), .A3(new_n331), .A4(new_n679), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n436), .B1(new_n435), .B2(new_n679), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n332), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n736), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n828), .B1(new_n735), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n735), .B2(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(new_n828), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n762), .A2(new_n812), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n203), .ZN(new_n843));
  INV_X1    g0643(.A(new_n762), .ZN(new_n844));
  INV_X1    g0644(.A(new_n789), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G87), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n775), .A2(G311), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n800), .A2(new_n304), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n793), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G303), .A2(new_n797), .B1(new_n849), .B2(G107), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n850), .B1(new_n591), .B2(new_n769), .C1(new_n475), .C2(new_n786), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(G116), .C2(new_n809), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G132), .A2(new_n775), .B1(new_n849), .B2(G50), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n218), .B2(new_n789), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n816), .B1(new_n217), .B2(new_n764), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G137), .A2(new_n797), .B1(new_n798), .B2(G143), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n254), .B2(new_n769), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G159), .B2(new_n809), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n854), .B(new_n855), .C1(new_n858), .C2(KEYINPUT34), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n858), .A2(KEYINPUT34), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n852), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n843), .B1(new_n844), .B2(new_n861), .C1(new_n837), .C2(new_n813), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n840), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n593), .B(new_n216), .C1(new_n536), .C2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n866), .A2(KEYINPUT102), .B1(new_n865), .B2(new_n536), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(KEYINPUT102), .B2(new_n866), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n703), .A2(G77), .A3(new_n391), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n344), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n259), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n412), .A2(new_n415), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n425), .A2(new_n426), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n678), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n431), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n412), .A2(new_n415), .A3(new_n430), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n427), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n879), .A4(new_n878), .ZN(new_n885));
  INV_X1    g0685(.A(new_n415), .ZN(new_n886));
  INV_X1    g0686(.A(new_n407), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT16), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n406), .A2(new_n218), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n408), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n249), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(KEYINPUT103), .A3(new_n249), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n876), .A2(new_n678), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n431), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n882), .A2(new_n885), .B1(new_n897), .B2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n678), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n428), .B2(new_n432), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n874), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n882), .A2(new_n885), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n678), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n895), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n634), .B2(new_n628), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n671), .A2(new_n837), .A3(new_n679), .ZN(new_n911));
  INV_X1    g0711(.A(new_n835), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n679), .A2(new_n348), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n384), .A2(new_n629), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n373), .B(KEYINPUT74), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n379), .A3(new_n382), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n914), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n910), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n634), .A2(new_n906), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n879), .B1(new_n884), .B2(new_n878), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n882), .B2(new_n885), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n878), .B1(new_n428), .B2(new_n432), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n874), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n909), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n902), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(new_n385), .A3(new_n679), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n438), .B1(new_n754), .B2(new_n738), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n638), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n902), .A2(new_n909), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n920), .A2(new_n732), .A3(new_n837), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n920), .A2(new_n732), .A3(new_n837), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(KEYINPUT40), .A3(new_n929), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n438), .A2(new_n732), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n948), .A2(new_n949), .A3(new_n685), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n939), .A2(new_n950), .B1(new_n259), .B2(new_n825), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n939), .A2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n873), .B1(new_n951), .B2(new_n952), .ZN(G367));
  INV_X1    g0753(.A(KEYINPUT109), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n695), .A2(new_n503), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n748), .B(new_n749), .C1(new_n517), .C2(new_n679), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n645), .A2(new_n660), .A3(new_n687), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(KEYINPUT108), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(new_n668), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n542), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n963), .B2(new_n679), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n687), .A2(new_n647), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n659), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n687), .A2(new_n647), .A3(new_n639), .ZN(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(new_n967), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n969), .B1(new_n964), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n693), .A2(new_n961), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n954), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n975), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n970), .A2(new_n973), .A3(KEYINPUT109), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(new_n975), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n701), .B(KEYINPUT41), .Z(new_n982));
  INV_X1    g0782(.A(new_n692), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n955), .B1(new_n983), .B2(new_n694), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(new_n686), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n757), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n696), .A2(new_n958), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT44), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n696), .A2(new_n958), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT110), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n988), .B1(KEYINPUT45), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n693), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n986), .B1(new_n995), .B2(KEYINPUT111), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n693), .A3(new_n993), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(new_n994), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n996), .B1(new_n999), .B2(KEYINPUT111), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n982), .B1(new_n1000), .B2(new_n757), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n981), .B1(new_n1001), .B2(new_n827), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n786), .A2(new_n254), .ZN(new_n1003));
  INV_X1    g0803(.A(G137), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1004), .A2(new_n774), .B1(new_n793), .B2(new_n217), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G143), .C2(new_n797), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n765), .A2(G68), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n789), .A2(new_n203), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n304), .B(new_n1008), .C1(G159), .C2(new_n770), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n809), .A2(G50), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT112), .B1(new_n849), .B2(G116), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT46), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n845), .A2(G97), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n774), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G303), .B2(new_n798), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1013), .B(new_n1017), .C1(new_n591), .C2(new_n782), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G311), .A2(new_n797), .B1(new_n770), .B2(G294), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n816), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n206), .C2(new_n764), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1011), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT47), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n762), .A3(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n814), .B(new_n762), .C1(new_n700), .C2(new_n566), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n239), .A2(new_n817), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n841), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n814), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1026), .B(new_n1029), .C1(new_n971), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1002), .A2(new_n1031), .ZN(G387));
  NAND2_X1  g0832(.A1(new_n983), .A2(new_n814), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n817), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n236), .B2(G45), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n699), .B2(new_n820), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n252), .A2(G50), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT50), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n466), .B1(new_n218), .B2(new_n203), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n699), .B(new_n1039), .C1(new_n1038), .C2(new_n1037), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(G107), .B2(new_n210), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n841), .B1(new_n1041), .B2(new_n815), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n765), .A2(new_n566), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n849), .A2(G77), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1043), .A2(new_n816), .A3(new_n1014), .A4(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n782), .A2(new_n218), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n254), .A2(new_n774), .B1(new_n786), .B2(new_n344), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n252), .A2(new_n769), .B1(new_n805), .B2(new_n791), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n765), .A2(G283), .B1(new_n849), .B2(G294), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n791), .A2(new_n787), .B1(new_n769), .B2(new_n783), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT113), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n581), .B2(new_n782), .C1(new_n1015), .C2(new_n786), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1020), .B1(new_n593), .B2(new_n789), .C1(new_n792), .C2(new_n774), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1056), .B2(KEYINPUT49), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1049), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1042), .B1(new_n844), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT114), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n985), .A2(new_n827), .B1(new_n1033), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n986), .A2(new_n701), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n985), .A2(new_n757), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(G393));
  OAI21_X1  g0866(.A(new_n986), .B1(new_n998), .B2(new_n994), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT111), .B1(new_n995), .B2(new_n997), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT111), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n757), .B(new_n985), .C1(new_n994), .C2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1067), .B(new_n701), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n961), .A2(new_n814), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n815), .B1(new_n205), .B2(new_n210), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1034), .A2(new_n243), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n828), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n787), .A2(new_n774), .B1(new_n769), .B2(new_n581), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n802), .B(new_n1076), .C1(G283), .C2(new_n849), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n277), .B1(G116), .B2(new_n765), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n475), .C2(new_n782), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n791), .A2(new_n1015), .B1(new_n786), .B2(new_n783), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  OAI22_X1  g0881(.A1(new_n791), .A2(new_n254), .B1(new_n786), .B2(new_n805), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n252), .B2(new_n782), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G143), .A2(new_n775), .B1(new_n849), .B2(G68), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G50), .A2(new_n770), .B1(new_n845), .B2(G87), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n765), .A2(G77), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n816), .A4(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1079), .A2(new_n1081), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1075), .B1(new_n1089), .B2(new_n762), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n999), .A2(new_n827), .B1(new_n1072), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1071), .A2(new_n1091), .ZN(G390));
  INV_X1    g0892(.A(KEYINPUT115), .ZN(new_n1093));
  AND4_X1   g0893(.A1(G330), .A2(new_n920), .A3(new_n732), .A4(new_n837), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n913), .A2(new_n920), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n385), .A2(new_n679), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n931), .A2(new_n932), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n383), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n915), .B1(new_n1098), .B2(new_n917), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n390), .B1(new_n918), .B2(new_n349), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n915), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n836), .A2(new_n332), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n753), .A2(new_n679), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1103), .B2(new_n912), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n929), .A2(new_n1096), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1093), .B(new_n1094), .C1(new_n1097), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n912), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n920), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n929), .A2(new_n1096), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n835), .B1(new_n736), .B2(new_n1102), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1096), .B1(new_n1101), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n932), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT39), .B1(new_n909), .B2(new_n928), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n727), .A2(new_n734), .A3(new_n837), .A4(new_n920), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1107), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1093), .B1(new_n1120), .B2(new_n1094), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n727), .A2(new_n734), .A3(new_n837), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1094), .B1(new_n1123), .B2(new_n1101), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1108), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n685), .B1(new_n730), .B2(new_n731), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n837), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1127), .B2(KEYINPUT116), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n920), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1124), .A2(new_n1112), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n438), .A2(new_n1127), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n335), .A2(new_n937), .A3(new_n1133), .A4(new_n637), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1132), .A2(KEYINPUT117), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT117), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1122), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n931), .A2(new_n932), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(new_n1113), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1094), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT115), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1107), .A3(new_n1118), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1132), .A2(KEYINPUT117), .A3(new_n1134), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1137), .A2(new_n1147), .A3(new_n701), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1141), .A2(new_n812), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n842), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n828), .B1(new_n1150), .B2(new_n251), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n786), .A2(new_n593), .B1(new_n769), .B2(new_n206), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n791), .A2(new_n591), .B1(new_n774), .B2(new_n475), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n809), .C2(G97), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n803), .B1(G68), .B2(new_n845), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1154), .A2(new_n304), .A3(new_n1087), .A4(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT118), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n849), .A2(G150), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT53), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G159), .B2(new_n765), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n809), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(G132), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n786), .A2(new_n1164), .B1(new_n769), .B2(new_n1004), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G125), .B2(new_n775), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n791), .A2(new_n1167), .B1(new_n789), .B2(new_n344), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n304), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1160), .A2(new_n1163), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1157), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT119), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(new_n844), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(KEYINPUT119), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1151), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1122), .A2(new_n827), .B1(new_n1149), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1148), .A2(new_n1176), .ZN(G378));
  NAND2_X1  g0977(.A1(new_n300), .A2(new_n335), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n265), .A2(new_n906), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n1181), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n812), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n828), .B1(new_n1150), .B2(G50), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n782), .A2(new_n323), .B1(new_n205), .B2(new_n769), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT121), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G116), .A2(new_n797), .B1(new_n798), .B2(G107), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n775), .A2(G283), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n1007), .A3(new_n1044), .A4(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n789), .A2(new_n217), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT120), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1020), .A2(new_n287), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1191), .A2(new_n1194), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1198), .B(new_n344), .C1(G33), .C2(G41), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G128), .A2(new_n798), .B1(new_n770), .B2(G132), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G125), .A2(new_n797), .B1(new_n849), .B2(new_n1162), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n254), .B2(new_n764), .C1(new_n1004), .C2(new_n782), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n845), .A2(G159), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n775), .C2(G124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1202), .B1(KEYINPUT58), .B2(new_n1199), .C1(new_n1207), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1189), .B1(new_n1212), .B2(new_n762), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1188), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n943), .A2(new_n945), .A3(G330), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1187), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1217), .A2(G330), .A3(new_n943), .A4(new_n945), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n936), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n936), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1214), .B1(new_n1223), .B2(new_n827), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1145), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1134), .ZN(new_n1226));
  OAI211_X1 g1026(.A(KEYINPUT57), .B(new_n1223), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n701), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n936), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n934), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n935), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1216), .A2(new_n1218), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1137), .B2(new_n1134), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT57), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1224), .B1(new_n1228), .B2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1132), .A2(new_n827), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1008), .B1(G283), .B2(new_n798), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n304), .A3(new_n1043), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n782), .A2(new_n206), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n791), .A2(new_n475), .B1(new_n769), .B2(new_n593), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n581), .A2(new_n774), .B1(new_n793), .B2(new_n205), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1167), .A2(new_n774), .B1(new_n793), .B2(new_n805), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1020), .B(new_n1244), .C1(G50), .C2(new_n765), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n1196), .C1(new_n254), .C2(new_n782), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n791), .A2(new_n1164), .B1(new_n786), .B2(new_n1004), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n770), .B2(new_n1162), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1243), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n828), .B1(G68), .B2(new_n1150), .C1(new_n1250), .C2(new_n844), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT123), .Z(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n813), .B2(new_n920), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1140), .A2(new_n1146), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n982), .B2(new_n1257), .ZN(G381));
  OR2_X1    g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  OR3_X1    g1059(.A1(G390), .A2(G384), .A3(new_n1259), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(G387), .A2(new_n1260), .A3(G381), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1224), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n701), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1234), .B2(KEYINPUT57), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT57), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1262), .B(G378), .C1(new_n1264), .C2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1261), .A2(new_n1268), .ZN(G407));
  INV_X1    g1069(.A(G343), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1261), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G213), .ZN(G409));
  NOR2_X1   g1072(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n701), .B1(new_n1273), .B2(KEYINPUT60), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1135), .A2(new_n1136), .A3(new_n1273), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(G384), .A3(new_n1255), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1274), .B1(new_n1257), .B2(KEYINPUT60), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1254), .A2(KEYINPUT124), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1237), .B2(new_n1253), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n863), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G213), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(G343), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(G2897), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1279), .A2(new_n1285), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1279), .B2(new_n1285), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1148), .A2(new_n1176), .A3(new_n1224), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n982), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1234), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1287), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1262), .B1(new_n1264), .B2(new_n1267), .ZN(new_n1296));
  INV_X1    g1096(.A(G378), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1265), .A2(new_n982), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1148), .A2(new_n1224), .A3(new_n1176), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n1300), .A2(new_n1301), .B1(new_n1286), .B2(G343), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(G378), .B2(G375), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1279), .A2(new_n1285), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1295), .B(new_n1305), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1299), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G393), .A2(G396), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1259), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1071), .B2(new_n1091), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1071), .A2(new_n1311), .A3(new_n1091), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1002), .A2(new_n1313), .A3(new_n1031), .A4(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n757), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1293), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n980), .B1(new_n1317), .B2(new_n826), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1031), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1314), .ZN(new_n1320));
  OAI22_X1  g1120(.A1(new_n1318), .A2(new_n1319), .B1(new_n1320), .B2(new_n1312), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1315), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1309), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1307), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1307), .A2(KEYINPUT125), .A3(new_n1324), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1322), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .A4(new_n1299), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1331), .B1(new_n1307), .B2(new_n1324), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1303), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1305), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1323), .B1(new_n1330), .B2(new_n1334), .ZN(G405));
  INV_X1    g1135(.A(new_n1305), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1297), .B1(new_n1337), .B2(new_n1224), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1336), .B1(new_n1338), .B2(new_n1268), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(G375), .A2(G378), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1341), .A3(new_n1305), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1339), .A2(new_n1322), .A3(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT127), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1339), .A2(new_n1322), .A3(new_n1342), .A4(KEYINPUT127), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1329), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1345), .A2(new_n1346), .A3(new_n1348), .ZN(G402));
endmodule


