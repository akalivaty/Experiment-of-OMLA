//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT80), .B(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(G101), .B1(new_n193), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT81), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n197), .A2(new_n199), .A3(new_n201), .A4(KEYINPUT82), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n194), .A2(new_n195), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n207), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT64), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n209), .B(new_n211), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT64), .A2(G143), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT64), .A2(G143), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n218), .A2(new_n219), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n208), .B1(new_n222), .B2(G146), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT81), .B(G107), .ZN(new_n225));
  OAI22_X1  g039(.A1(G104), .A2(new_n225), .B1(new_n193), .B2(G107), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT84), .B1(new_n226), .B2(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n196), .A2(KEYINPUT80), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT80), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G104), .ZN(new_n230));
  AOI21_X1  g044(.A(G107), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(G104), .B1(new_n199), .B2(new_n201), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT84), .B(G101), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n206), .B(new_n224), .C1(new_n227), .C2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n193), .A2(G107), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n194), .A2(new_n204), .A3(new_n238), .A4(new_n205), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(G146), .B1(new_n213), .B2(new_n214), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT65), .B1(new_n216), .B2(G143), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n243), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n209), .B(new_n244), .C1(new_n215), .C2(new_n216), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G101), .ZN(new_n252));
  OR2_X1    g066(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n239), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n241), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT11), .B1(new_n258), .B2(G137), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(G137), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT66), .A2(G131), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT66), .A2(G131), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n263), .B2(new_n264), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n272));
  OAI21_X1  g086(.A(G128), .B1(new_n208), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n243), .C1(new_n247), .C2(new_n248), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n217), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(KEYINPUT10), .ZN(new_n276));
  OAI21_X1  g090(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n233), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n206), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n237), .A2(new_n257), .A3(new_n271), .A4(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT86), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n205), .B1(new_n231), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT82), .B1(new_n225), .B2(new_n197), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n279), .A2(new_n233), .B1(new_n288), .B2(new_n195), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n235), .A2(new_n236), .B1(new_n289), .B2(new_n276), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(KEYINPUT86), .A3(new_n271), .A4(new_n257), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G227), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G953), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n235), .B1(new_n289), .B2(new_n275), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n259), .A2(new_n262), .B1(new_n258), .B2(G137), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n269), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT12), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(KEYINPUT12), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n292), .A2(KEYINPUT87), .A3(new_n297), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n300), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n290), .A2(new_n257), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n304), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n292), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n296), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n192), .B1(new_n316), .B2(new_n190), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n292), .A2(new_n313), .A3(new_n297), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n292), .A2(new_n309), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(new_n297), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(new_n190), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n189), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(G125), .A2(G140), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT74), .B(G125), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n324), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n216), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(KEYINPUT16), .B2(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n210), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT24), .B(G110), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n334), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(G110), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n332), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G110), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(new_n341), .A3(new_n345), .A4(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G125), .B(G140), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT76), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G146), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n331), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G137), .ZN(new_n356));
  INV_X1    g170(.A(G953), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(G221), .A3(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n344), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n353), .B1(new_n330), .B2(G146), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n332), .A2(new_n343), .B1(new_n361), .B2(new_n350), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n359), .B(KEYINPUT77), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n360), .B(new_n191), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n344), .A2(new_n355), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n363), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n360), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(KEYINPUT78), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G234), .B2(new_n191), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n374), .A3(new_n366), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n369), .A2(new_n360), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n373), .A2(G902), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(G472), .A2(G902), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n357), .A3(G210), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT27), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT26), .B(G101), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n304), .A2(new_n249), .A3(new_n250), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n264), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n258), .A2(KEYINPUT68), .A3(G137), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n261), .A2(G134), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(G131), .A2(new_n394), .B1(new_n303), .B2(new_n267), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n275), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n333), .A2(G116), .ZN(new_n398));
  INV_X1    g212(.A(G116), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G119), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT2), .B(G113), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT69), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT69), .B1(new_n401), .B2(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n401), .A2(new_n403), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n388), .B1(new_n397), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n413));
  INV_X1    g227(.A(KEYINPUT67), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n271), .B2(new_n251), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n304), .A2(KEYINPUT67), .A3(new_n249), .A4(new_n250), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT30), .B1(new_n417), .B2(new_n396), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n389), .A2(new_n396), .A3(KEYINPUT30), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n410), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n412), .B(new_n413), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT71), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n415), .A2(new_n416), .B1(new_n275), .B2(new_n395), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n410), .B(new_n419), .C1(new_n423), .C2(KEYINPUT30), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT71), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n412), .A4(new_n413), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n412), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n397), .B2(new_n411), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n389), .A2(new_n396), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n431), .A2(KEYINPUT28), .A3(new_n410), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n430), .A2(new_n432), .B1(new_n423), .B2(new_n411), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n428), .A2(KEYINPUT31), .B1(new_n433), .B2(new_n388), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n427), .B2(new_n434), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT32), .B(new_n382), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n430), .A2(new_n432), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n410), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n388), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(G902), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n397), .A2(new_n411), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n424), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n387), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n443), .B1(new_n433), .B2(new_n388), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G472), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n438), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n382), .B1(new_n436), .B2(new_n437), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n381), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n274), .A2(new_n217), .A3(new_n324), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n324), .B1(new_n249), .B2(new_n250), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n459), .A2(new_n460), .ZN(new_n464));
  INV_X1    g278(.A(G224), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G953), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT90), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n409), .A2(new_n408), .B1(new_n239), .B2(new_n255), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n241), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(G113), .C1(KEYINPUT5), .C2(new_n398), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n280), .A2(new_n408), .A3(new_n206), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n473), .B2(new_n476), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n471), .B(new_n482), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n206), .B1(new_n227), .B2(new_n234), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n475), .A2(new_n408), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n476), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n478), .B(KEYINPUT8), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n494), .A2(new_n481), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT7), .B1(new_n465), .B2(G953), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n464), .B(new_n496), .C1(new_n462), .C2(new_n461), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n488), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G210), .B1(G237), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n488), .A2(new_n501), .A3(new_n503), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(KEYINPUT91), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G214), .B1(G237), .B2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n506), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n383), .A2(new_n357), .A3(G143), .A4(G214), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n383), .A2(new_n357), .A3(G214), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n215), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n267), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(KEYINPUT19), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n352), .B2(KEYINPUT19), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n331), .B(new_n520), .C1(G146), .C2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n326), .A2(new_n216), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n516), .A2(new_n525), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n353), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G113), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n196), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  INV_X1    g348(.A(new_n519), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(KEYINPUT17), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n519), .A2(KEYINPUT92), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n518), .A2(new_n537), .A3(new_n519), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n329), .A3(new_n331), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n531), .B(new_n528), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n513), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n513), .A3(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n528), .B1(new_n539), .B2(new_n541), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n532), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n542), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n191), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n546), .A2(new_n547), .B1(G475), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(G234), .A2(G237), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(G952), .A3(new_n357), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT21), .B(G898), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(G902), .A3(G953), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT97), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n213), .A2(G128), .A3(new_n214), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n560), .B(new_n258), .C1(G128), .C2(new_n207), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT93), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(KEYINPUT13), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(new_n258), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n560), .B(KEYINPUT13), .C1(G128), .C2(new_n207), .ZN(new_n565));
  XNOR2_X1  g379(.A(G116), .B(G122), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n225), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n225), .A2(new_n566), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n564), .A2(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G122), .ZN(new_n571));
  OR3_X1    g385(.A1(new_n571), .A2(KEYINPUT14), .A3(G116), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT95), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(G116), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT14), .B1(new_n571), .B2(G116), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n572), .A2(KEYINPUT95), .ZN(new_n577));
  OAI21_X1  g391(.A(G107), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n568), .B(KEYINPUT94), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n560), .B1(G128), .B2(new_n207), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G134), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n561), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n187), .A2(new_n372), .A3(G953), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n570), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n570), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n191), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G478), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT15), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n570), .A2(new_n583), .ZN(new_n593));
  INV_X1    g407(.A(new_n584), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n570), .A2(new_n583), .A3(new_n584), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(KEYINPUT96), .A3(new_n191), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n598), .A3(new_n589), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n552), .A2(new_n559), .A3(new_n590), .A4(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n512), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n322), .A2(new_n458), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT98), .B(G101), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  INV_X1    g418(.A(new_n381), .ZN(new_n605));
  INV_X1    g419(.A(new_n382), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n427), .A2(new_n434), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT72), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n191), .B1(new_n436), .B2(new_n437), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n610), .B1(G472), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n322), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n508), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n505), .B2(new_n506), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n592), .A2(new_n598), .A3(new_n588), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n191), .A2(G478), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n595), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n597), .A2(new_n619), .A3(KEYINPUT33), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n595), .B(new_n596), .C1(new_n618), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n552), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n615), .A2(new_n559), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n196), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND2_X1  g445(.A1(new_n599), .A2(new_n590), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n552), .A2(new_n615), .A3(new_n559), .A4(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n613), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n611), .A2(G472), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n368), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n379), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n376), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n638), .A2(new_n454), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n322), .A2(new_n644), .A3(new_n601), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  NAND2_X1  g461(.A1(new_n552), .A2(new_n632), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n557), .A2(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n554), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n438), .A2(new_n452), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n608), .A2(new_n609), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n455), .B1(new_n654), .B2(new_n382), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n642), .B(new_n652), .C1(new_n653), .C2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n310), .A2(new_n309), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT87), .B1(new_n292), .B2(new_n297), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n315), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n190), .A3(new_n191), .ZN(new_n660));
  INV_X1    g474(.A(new_n192), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n321), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n188), .A3(new_n615), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n210), .ZN(G30));
  XNOR2_X1  g479(.A(new_n650), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n322), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n446), .A2(new_n388), .A3(new_n440), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n447), .B2(new_n387), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n191), .B1(new_n672), .B2(new_n673), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n438), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n670), .B1(new_n677), .B2(new_n655), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n457), .A2(KEYINPUT102), .A3(new_n438), .A4(new_n676), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n503), .B1(new_n488), .B2(new_n501), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n509), .A2(new_n681), .A3(new_n510), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n506), .A2(KEYINPUT91), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT38), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n507), .A2(new_n685), .A3(new_n511), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n543), .A2(new_n513), .A3(new_n544), .ZN(new_n688));
  INV_X1    g502(.A(G475), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n549), .B2(new_n542), .ZN(new_n690));
  OAI22_X1  g504(.A1(new_n688), .A2(new_n545), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n376), .A2(new_n691), .A3(new_n632), .A4(new_n641), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n687), .A2(new_n614), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n668), .A2(new_n669), .A3(new_n680), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n215), .ZN(G45));
  AND3_X1   g514(.A1(new_n662), .A2(new_n188), .A3(new_n615), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n624), .A2(new_n552), .A3(new_n651), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n642), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n453), .B2(new_n457), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NAND2_X1  g520(.A1(new_n660), .A2(new_n188), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT104), .B1(new_n316), .B2(new_n190), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n659), .A2(new_n191), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(G469), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n707), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n458), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n627), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n634), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n399), .ZN(G18));
  INV_X1    g532(.A(new_n642), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n453), .B2(new_n457), .ZN(new_n720));
  INV_X1    g534(.A(new_n600), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n712), .A3(new_n721), .A4(new_n615), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AND2_X1   g537(.A1(new_n691), .A2(new_n632), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n615), .A2(new_n559), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n428), .A2(KEYINPUT31), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n427), .B(new_n726), .C1(new_n387), .C2(new_n442), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n382), .B(KEYINPUT105), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n638), .A2(new_n605), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n611), .A2(G472), .B1(new_n727), .B2(new_n728), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT106), .B1(new_n733), .B2(new_n605), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n712), .B(new_n725), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AOI21_X1  g550(.A(new_n189), .B1(new_n316), .B2(new_n190), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n710), .B1(new_n709), .B2(G469), .ZN(new_n738));
  AOI211_X1 g552(.A(KEYINPUT104), .B(new_n190), .C1(new_n659), .C2(new_n191), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n615), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n733), .A2(new_n642), .A3(new_n702), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(G125), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n188), .B(new_n508), .C1(new_n682), .C2(new_n683), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n292), .A2(new_n313), .A3(new_n297), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n297), .B1(new_n292), .B2(new_n309), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT108), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(G469), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT109), .A4(G469), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n746), .B1(new_n317), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n610), .A2(KEYINPUT32), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n605), .B(new_n702), .C1(new_n757), .C2(new_n653), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n745), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n317), .ZN(new_n761));
  INV_X1    g575(.A(new_n746), .ZN(new_n762));
  INV_X1    g576(.A(new_n702), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(KEYINPUT42), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n458), .A2(new_n761), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND4_X1  g581(.A1(new_n458), .A2(new_n761), .A3(new_n762), .A4(new_n652), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  AOI21_X1  g583(.A(new_n614), .B1(new_n507), .B2(new_n511), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n616), .A2(new_n623), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n552), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n552), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n642), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n612), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n771), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(KEYINPUT44), .B2(new_n781), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT45), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n190), .B1(new_n320), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n192), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n660), .B1(new_n787), .B2(KEYINPUT46), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n789), .B(new_n192), .C1(new_n784), .C2(new_n786), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n188), .B(new_n666), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n261), .ZN(G39));
  NAND2_X1  g607(.A1(new_n453), .A2(new_n457), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n770), .A2(new_n381), .A3(new_n702), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n188), .B1(new_n788), .B2(new_n790), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(KEYINPUT47), .B(new_n188), .C1(new_n788), .C2(new_n790), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n794), .B(new_n795), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n325), .ZN(G42));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n692), .A2(new_n615), .A3(new_n188), .A4(new_n650), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n755), .B2(new_n317), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n680), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n705), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  OAI22_X1  g621(.A1(new_n740), .A2(new_n741), .B1(new_n656), .B2(new_n663), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n808), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n680), .A2(new_n804), .B1(new_n701), .B2(new_n704), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n624), .B2(new_n552), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n691), .B(KEYINPUT112), .C1(new_n616), .C2(new_n623), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n648), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n559), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n512), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n322), .A3(new_n605), .A4(new_n612), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n735), .A2(new_n820), .A3(new_n722), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n322), .B(new_n601), .C1(new_n458), .C2(new_n644), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n458), .B(new_n712), .C1(new_n626), .C2(new_n633), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n719), .A2(new_n691), .A3(new_n632), .A4(new_n651), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n322), .A2(new_n794), .A3(new_n770), .A4(new_n825), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n638), .A2(new_n642), .A3(new_n702), .A4(new_n729), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n761), .A3(new_n762), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n768), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n821), .A2(new_n766), .A3(new_n824), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n802), .B1(new_n813), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n807), .B1(new_n806), .B2(new_n808), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n810), .A2(KEYINPUT52), .A3(new_n811), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n735), .A2(new_n820), .A3(new_n722), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n822), .A2(new_n823), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n768), .A2(new_n826), .A3(new_n828), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n760), .A3(new_n765), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n831), .A2(new_n832), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT114), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n831), .A2(new_n844), .A3(new_n841), .A4(new_n832), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n831), .A2(new_n841), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n832), .B1(new_n831), .B2(new_n841), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n773), .A2(new_n774), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n554), .B1(new_n855), .B2(new_n778), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n732), .B2(new_n734), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n508), .B1(new_n684), .B2(new_n686), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n712), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n854), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n856), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n730), .A2(new_n731), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n605), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(KEYINPUT50), .A3(new_n712), .A4(new_n858), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n712), .A2(new_n770), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n680), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n381), .A2(new_n554), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n772), .A2(new_n691), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n712), .A2(new_n770), .A3(new_n856), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n733), .A2(new_n642), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT117), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n712), .A2(new_n770), .A3(new_n856), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(new_n875), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n873), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n853), .B1(new_n867), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n798), .A2(new_n799), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n708), .A2(new_n711), .B1(new_n190), .B2(new_n316), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n189), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT119), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n857), .B2(new_n771), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n864), .A2(KEYINPUT115), .A3(new_n770), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n798), .A2(new_n892), .A3(new_n799), .A4(new_n885), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n874), .A2(KEYINPUT117), .A3(new_n876), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n879), .B1(new_n878), .B2(new_n875), .ZN(new_n896));
  INV_X1    g710(.A(new_n871), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n868), .A2(new_n680), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n895), .A2(new_n896), .B1(new_n898), .B2(new_n872), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(KEYINPUT118), .A3(new_n866), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n882), .A2(new_n894), .A3(KEYINPUT51), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT51), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n889), .A2(new_n890), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n886), .B1(new_n883), .B2(KEYINPUT116), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT116), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n798), .A2(new_n905), .A3(new_n799), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n899), .A2(new_n866), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n902), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n605), .B1(new_n757), .B2(new_n653), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n878), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT48), .Z(new_n912));
  NOR2_X1   g726(.A1(new_n857), .A2(new_n740), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT120), .ZN(new_n914));
  INV_X1    g728(.A(G952), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n915), .B(G953), .C1(new_n898), .C2(new_n625), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n912), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n901), .A2(new_n909), .A3(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n846), .A2(new_n849), .A3(new_n852), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n850), .B(KEYINPUT113), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n922), .A3(new_n846), .A4(new_n918), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n357), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n773), .A2(new_n381), .A3(new_n189), .A4(new_n614), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT49), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n884), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT111), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n884), .A2(new_n927), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n929), .A2(new_n870), .A3(new_n687), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n925), .A2(new_n931), .ZN(G75));
  INV_X1    g746(.A(new_n847), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n191), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(new_n471), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT55), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(KEYINPUT56), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n935), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n935), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n357), .A2(G952), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G51));
  XNOR2_X1  g759(.A(new_n192), .B(KEYINPUT57), .ZN(new_n946));
  INV_X1    g760(.A(new_n842), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n850), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT123), .B(new_n946), .C1(new_n947), .C2(new_n850), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n659), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n934), .A2(new_n784), .A3(new_n786), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n944), .B1(new_n952), .B2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  INV_X1    g769(.A(new_n543), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n944), .ZN(G60));
  NAND2_X1  g773(.A1(new_n620), .A2(new_n622), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n921), .A2(new_n846), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT59), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n960), .B(new_n963), .C1(new_n947), .C2(new_n850), .ZN(new_n965));
  INV_X1    g779(.A(new_n944), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n964), .A2(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n933), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n640), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n377), .B(KEYINPUT124), .Z(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n933), .B2(new_n970), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n966), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n555), .B2(new_n465), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n838), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n936), .B1(G898), .B2(new_n357), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  OAI21_X1  g795(.A(new_n419), .B1(new_n423), .B2(KEYINPUT30), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n522), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n808), .B1(new_n701), .B2(new_n704), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n697), .A2(new_n698), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n458), .A2(new_n770), .A3(new_n817), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(new_n667), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n792), .A2(new_n800), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n983), .B1(new_n991), .B2(new_n357), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n357), .B1(G227), .B2(G900), .ZN(new_n993));
  INV_X1    g807(.A(G900), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n983), .B1(new_n994), .B2(new_n357), .ZN(new_n995));
  INV_X1    g809(.A(new_n792), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n996), .A2(new_n984), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n615), .A2(new_n724), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n791), .A2(new_n998), .A3(new_n910), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n766), .A2(new_n768), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n800), .A2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n995), .B1(new_n1002), .B2(new_n357), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n992), .A2(new_n993), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n993), .B1(new_n992), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(new_n447), .A2(new_n387), .ZN(new_n1007));
  XNOR2_X1  g821(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n448), .A2(new_n388), .ZN(new_n1012));
  AND4_X1   g826(.A1(new_n1007), .A2(new_n847), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n986), .A2(new_n838), .A3(new_n987), .A4(new_n990), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1010), .B(KEYINPUT126), .Z(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1007), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n997), .A2(new_n838), .A3(new_n999), .A4(new_n1001), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1012), .B1(new_n1018), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT127), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n944), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n1019), .B2(new_n944), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1013), .B(new_n1017), .C1(new_n1021), .C2(new_n1022), .ZN(G57));
endmodule


