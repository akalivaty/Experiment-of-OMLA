//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1306, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n214), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n223), .A2(G1), .A3(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n212), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n203), .A2(G50), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n220), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n217), .B(new_n230), .C1(KEYINPUT1), .C2(new_n215), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G107), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G238), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n249), .B1(new_n250), .B2(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n225), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  INV_X1    g0057(.A(new_n221), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(new_n254), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(G244), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G179), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n222), .A2(new_n224), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT66), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n222), .A2(new_n224), .A3(new_n275), .A4(new_n272), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G13), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT69), .A3(G20), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n274), .A2(new_n276), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n212), .A2(G1), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n279), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n283), .A2(new_n286), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT15), .B(G87), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n212), .A2(G33), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XOR2_X1   g0094(.A(KEYINPUT8), .B(G58), .Z(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(new_n296), .B1(G20), .B2(G77), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n274), .A2(new_n276), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n290), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n271), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n295), .ZN(new_n309));
  INV_X1    g0109(.A(G150), .ZN(new_n310));
  INV_X1    g0110(.A(new_n296), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n309), .A2(new_n293), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n203), .A2(G50), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n212), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n300), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n277), .ZN(new_n316));
  INV_X1    g0116(.A(G50), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n274), .A2(new_n276), .ZN(new_n320));
  INV_X1    g0120(.A(new_n284), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(G50), .A3(new_n277), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n325));
  INV_X1    g0125(.A(G223), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n285), .B2(new_n247), .C1(new_n251), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n255), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n263), .B1(G226), .B2(new_n266), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G179), .ZN(new_n331));
  AOI21_X1  g0131(.A(G169), .B1(new_n328), .B2(new_n329), .ZN(new_n332));
  OR3_X1    g0132(.A1(new_n324), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n256), .A2(G190), .A3(new_n267), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n268), .A2(G200), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n306), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n308), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(G232), .A4(G1698), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n339), .A2(new_n341), .A3(G226), .A4(new_n248), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n345), .A2(new_n255), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n264), .A2(G274), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT70), .B1(new_n347), .B2(new_n260), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n261), .A2(new_n264), .A3(new_n349), .A4(G274), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n264), .A2(G238), .A3(new_n260), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT13), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n255), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(new_n348), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT14), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n353), .A2(G179), .A3(new_n357), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n362), .A3(G169), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n320), .A2(G68), .A3(new_n321), .A4(new_n287), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n202), .A2(G20), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n366), .B1(new_n293), .B2(new_n285), .C1(new_n311), .C2(new_n317), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(new_n274), .A3(new_n276), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT12), .B1(new_n287), .B2(G68), .ZN(new_n371));
  OR4_X1    g0171(.A1(KEYINPUT12), .A2(new_n366), .A3(G1), .A4(new_n280), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n367), .A2(new_n274), .A3(KEYINPUT11), .A4(new_n276), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n365), .A2(new_n370), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n369), .A2(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n378), .A2(KEYINPUT72), .A3(new_n374), .A4(new_n365), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n364), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n353), .A2(G190), .A3(new_n357), .ZN(new_n383));
  AND4_X1   g0183(.A1(new_n370), .A2(new_n365), .A3(new_n373), .A4(new_n374), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n353), .B2(new_n357), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n382), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n358), .A2(G200), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n389), .A2(KEYINPUT71), .A3(new_n384), .A4(new_n383), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT9), .B1(new_n319), .B2(new_n323), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT9), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n315), .A2(new_n393), .A3(new_n322), .A4(new_n318), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n330), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n386), .B1(new_n328), .B2(new_n329), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n337), .A2(new_n381), .A3(new_n391), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n263), .B1(G232), .B2(new_n266), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n247), .A2(G226), .A3(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n247), .A2(G223), .A3(new_n248), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n407), .B(new_n408), .C1(new_n338), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n255), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n411), .A3(new_n396), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n266), .A2(G232), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n262), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n255), .B2(new_n410), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n412), .B1(new_n415), .B2(G200), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n309), .A2(new_n284), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n320), .A2(new_n417), .A3(new_n277), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n277), .B2(new_n295), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n247), .B2(G20), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n340), .A2(G33), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n424));
  OAI211_X1 g0224(.A(KEYINPUT7), .B(new_n212), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT75), .B1(new_n426), .B2(G68), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n428), .B(new_n202), .C1(new_n422), .C2(new_n425), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G58), .A2(G68), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n203), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G20), .ZN(new_n436));
  INV_X1    g0236(.A(G159), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n437), .A2(G20), .A3(G33), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT74), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT74), .ZN(new_n441));
  AOI211_X1 g0241(.A(new_n441), .B(new_n438), .C1(new_n435), .C2(G20), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT16), .B1(new_n430), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT73), .B1(G58), .B2(G68), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n212), .B1(new_n447), .B2(new_n203), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n441), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n339), .A2(new_n341), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT7), .B1(new_n450), .B2(new_n212), .ZN(new_n451));
  AOI211_X1 g0251(.A(new_n421), .B(G20), .C1(new_n339), .C2(new_n341), .ZN(new_n452));
  OAI21_X1  g0252(.A(G68), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n436), .A2(KEYINPUT74), .A3(new_n439), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n449), .A2(new_n453), .A3(KEYINPUT16), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n300), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n416), .B(new_n420), .C1(new_n444), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n428), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n426), .A2(KEYINPUT75), .A3(G68), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n443), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT16), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n455), .A2(new_n300), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n419), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(KEYINPUT17), .A3(new_n416), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n415), .A2(G179), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n406), .A2(new_n411), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G169), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n456), .B1(new_n463), .B2(new_n462), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT18), .B(new_n473), .C1(new_n474), .C2(new_n419), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT76), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n420), .B1(new_n444), .B2(new_n456), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(KEYINPUT76), .A3(KEYINPUT18), .A4(new_n473), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT18), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n470), .A2(new_n472), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n466), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n469), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n405), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n339), .A2(new_n341), .A3(G264), .A4(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(new_n248), .ZN(new_n488));
  INV_X1    g0288(.A(G303), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n247), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n255), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n211), .A2(G45), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n259), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n265), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G270), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G169), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  INV_X1    g0301(.A(G179), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT85), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n338), .A2(G1), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n320), .A2(new_n287), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT84), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n283), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G20), .B1(G33), .B2(G283), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n338), .A2(G97), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n513), .A2(new_n514), .B1(G20), .B2(new_n506), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n515), .A2(new_n273), .A3(KEYINPUT20), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT20), .B1(new_n515), .B2(new_n273), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n516), .A2(new_n517), .B1(G116), .B2(new_n287), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n504), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  AOI211_X1 g0320(.A(KEYINPUT85), .B(new_n518), .C1(new_n509), .C2(new_n511), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n503), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND4_X1   g0322(.A1(new_n510), .A2(new_n320), .A3(new_n287), .A4(new_n507), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n510), .B1(new_n283), .B2(new_n507), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT85), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n512), .A2(new_n504), .A3(new_n519), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n499), .A2(G200), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n499), .A2(new_n396), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n500), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n522), .B(new_n530), .C1(new_n531), .C2(KEYINPUT21), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n339), .A2(new_n341), .A3(G238), .A4(new_n248), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n255), .ZN(new_n537));
  INV_X1    g0337(.A(G45), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G1), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n264), .A2(G274), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n264), .A2(G250), .A3(new_n492), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(G190), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n542), .B1(new_n255), .B2(new_n536), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n386), .ZN(new_n546));
  INV_X1    g0346(.A(new_n505), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n320), .A2(G87), .A3(new_n277), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n409), .A2(new_n549), .A3(new_n250), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT81), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n552), .A2(new_n409), .A3(new_n549), .A4(new_n250), .ZN(new_n553));
  NAND3_X1  g0353(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n551), .A2(new_n553), .B1(new_n212), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n339), .A2(new_n341), .A3(new_n212), .A4(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n293), .B2(new_n549), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n274), .B(new_n276), .C1(new_n555), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n288), .A2(new_n291), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n548), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n546), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n537), .A2(G179), .A3(new_n543), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n545), .B2(new_n269), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n560), .A2(new_n561), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n291), .B(KEYINPUT82), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n320), .A2(new_n567), .A3(new_n277), .A4(new_n547), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n565), .A2(KEYINPUT80), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT80), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n564), .B(new_n570), .C1(new_n269), .C2(new_n545), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n563), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(new_n248), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G283), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n255), .ZN(new_n580));
  AND2_X1   g0380(.A1(KEYINPUT5), .A2(G41), .ZN(new_n581));
  NOR2_X1   g0381(.A1(KEYINPUT5), .A2(G41), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n539), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(G257), .A3(new_n264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n496), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT79), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n585), .B1(new_n579), .B2(new_n255), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT79), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(G190), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n316), .A2(new_n549), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n296), .A2(G77), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n597), .A2(new_n549), .A3(G107), .ZN(new_n598));
  XNOR2_X1  g0398(.A(G97), .B(G107), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n596), .B1(new_n600), .B2(new_n212), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n250), .B1(new_n422), .B2(new_n425), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n300), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT77), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n595), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(KEYINPUT77), .B(new_n300), .C1(new_n601), .C2(new_n602), .ZN(new_n606));
  AOI211_X1 g0406(.A(new_n316), .B(new_n505), .C1(new_n274), .C2(new_n276), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G97), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n592), .A2(new_n593), .A3(new_n605), .A4(new_n609), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n588), .B(new_n585), .C1(new_n255), .C2(new_n579), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT79), .B1(new_n580), .B2(new_n586), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n269), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n603), .A2(new_n604), .ZN(new_n614));
  INV_X1    g0414(.A(new_n595), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n606), .A4(new_n608), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n587), .A2(G179), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n572), .A2(new_n610), .A3(new_n619), .A4(KEYINPUT83), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n339), .A2(new_n341), .A3(new_n212), .A4(G87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT22), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT22), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n247), .A2(new_n623), .A3(new_n212), .A4(G87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT24), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n535), .A2(G20), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT23), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n212), .B2(G107), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n250), .A2(KEYINPUT23), .A3(G20), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n626), .B1(new_n625), .B2(new_n631), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n300), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n316), .A2(new_n250), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT25), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n607), .B2(G107), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n497), .A2(G264), .B1(new_n259), .B2(new_n495), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(G1698), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n339), .A2(new_n341), .A3(G250), .A4(new_n248), .ZN(new_n641));
  NAND2_X1  g0441(.A1(G33), .A2(G294), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n255), .ZN(new_n644));
  AOI21_X1  g0444(.A(G169), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n497), .A2(G264), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n644), .A2(new_n646), .A3(new_n496), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n502), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n638), .A2(new_n648), .A3(KEYINPUT86), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT86), .B1(new_n638), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(G190), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n639), .A2(new_n644), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G200), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n634), .A2(new_n651), .A3(new_n637), .A4(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n649), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n620), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n572), .A2(new_n610), .A3(new_n619), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT83), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n486), .A2(new_n532), .A3(new_n661), .ZN(G372));
  INV_X1    g0462(.A(new_n333), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n404), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n401), .A2(new_n403), .A3(KEYINPUT87), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n482), .A2(new_n475), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n389), .A2(new_n384), .A3(new_n383), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n364), .A2(new_n380), .B1(new_n307), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n670), .B2(new_n468), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n663), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n386), .B1(new_n537), .B2(new_n543), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(G190), .B2(new_n545), .ZN(new_n674));
  INV_X1    g0474(.A(new_n562), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n568), .A2(new_n560), .A3(new_n561), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n674), .A2(new_n675), .B1(new_n565), .B2(new_n676), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n610), .A2(new_n619), .A3(new_n654), .A4(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n522), .B1(new_n531), .B2(KEYINPUT21), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n638), .A2(new_n648), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n572), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n617), .B1(new_n609), .B2(new_n605), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n677), .A3(new_n683), .A4(new_n613), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n565), .A2(new_n676), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n672), .B1(new_n486), .B2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(G213), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n280), .A2(G1), .A3(G20), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT27), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n697), .B2(new_n696), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n526), .B2(new_n527), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n532), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n500), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n520), .B2(new_n521), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n526), .A2(new_n527), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n707), .A2(new_n501), .B1(new_n708), .B2(new_n503), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(KEYINPUT89), .A3(new_n530), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n705), .A2(new_n710), .B1(new_n709), .B2(new_n703), .ZN(new_n711));
  XOR2_X1   g0511(.A(KEYINPUT90), .B(G330), .Z(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n656), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n638), .A2(new_n701), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n716), .A2(new_n717), .B1(new_n680), .B2(new_n702), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n681), .A2(new_n702), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n679), .A2(new_n702), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n656), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n218), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n551), .A2(new_n506), .A3(new_n553), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(G1), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n229), .B2(new_n727), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n532), .A2(new_n701), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n657), .A2(new_n733), .A3(new_n660), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n639), .A2(new_n491), .A3(new_n498), .A4(new_n644), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n564), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n589), .A3(new_n591), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n611), .A2(new_n612), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n736), .ZN(new_n741));
  AOI21_X1  g0541(.A(G179), .B1(new_n537), .B2(new_n543), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n499), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT91), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n587), .A2(new_n746), .A3(new_n652), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT92), .B1(new_n647), .B2(new_n590), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n499), .A2(new_n742), .A3(KEYINPUT91), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n745), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n739), .A2(new_n741), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n751), .B2(new_n701), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT93), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT30), .B1(new_n740), .B2(new_n736), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n739), .A2(KEYINPUT93), .A3(new_n750), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n741), .A3(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n701), .A2(KEYINPUT31), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n752), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n712), .B1(new_n734), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT29), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n649), .A2(new_n650), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n678), .B1(new_n679), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n684), .A2(new_n683), .A3(new_n572), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n674), .A2(new_n675), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n688), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT26), .B1(new_n619), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n765), .A2(new_n768), .A3(new_n688), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n762), .B1(new_n770), .B2(new_n702), .ZN(new_n771));
  AOI211_X1 g0571(.A(KEYINPUT29), .B(new_n701), .C1(new_n682), .C2(new_n690), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n761), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n732), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(new_n280), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n211), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n726), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n715), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n711), .A2(new_n713), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n711), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n218), .A2(new_n247), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n218), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n218), .A2(new_n450), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n229), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n538), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n242), .A2(new_n538), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n226), .B1(G20), .B2(new_n269), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n784), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n778), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n797), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n396), .A2(G179), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n212), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n212), .A2(new_n502), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(KEYINPUT33), .A2(G317), .ZN(new_n810));
  NAND2_X1  g0610(.A1(KEYINPUT33), .A2(G317), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n807), .A2(new_n396), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n805), .B(new_n812), .C1(G326), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n212), .A2(G190), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(new_n502), .A3(new_n386), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(new_n806), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n819), .A2(G190), .A3(G200), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n819), .A2(new_n396), .A3(G200), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n247), .B(new_n823), .C1(G322), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT96), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n386), .B2(G179), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n502), .A2(KEYINPUT96), .A3(G200), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n827), .A2(new_n828), .A3(new_n815), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G283), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n212), .A2(new_n396), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n827), .A2(new_n832), .A3(new_n828), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G303), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n814), .A2(new_n825), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n824), .B(KEYINPUT95), .Z(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G58), .B1(G107), .B2(new_n830), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n816), .A2(new_n437), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT32), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n450), .B1(new_n820), .B2(G77), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n834), .A2(G87), .ZN(new_n842));
  INV_X1    g0642(.A(new_n803), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G97), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G50), .A2(new_n813), .B1(new_n808), .B2(G68), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n838), .A2(new_n840), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n801), .B1(new_n836), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n800), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n779), .A2(new_n781), .B1(new_n786), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  NOR3_X1   g0651(.A1(new_n271), .A2(new_n306), .A3(new_n701), .ZN(new_n852));
  INV_X1    g0652(.A(new_n305), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n289), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n701), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n336), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n852), .B1(new_n857), .B2(new_n308), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n692), .B2(new_n701), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n610), .A2(new_n619), .A3(new_n654), .A4(new_n677), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n709), .B2(new_n680), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n571), .A3(new_n676), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n766), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT26), .B1(new_n865), .B2(new_n619), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n688), .A3(new_n687), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n702), .B(new_n858), .C1(new_n862), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n860), .A2(new_n761), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n869), .B(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n778), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n860), .A2(new_n868), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n871), .B(new_n872), .C1(new_n761), .C2(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n820), .A2(G159), .B1(new_n813), .B2(G137), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n310), .B2(new_n809), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT99), .B(G143), .Z(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n837), .B2(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT34), .Z(new_n880));
  AOI21_X1  g0680(.A(new_n450), .B1(new_n817), .B2(G132), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n830), .A2(G68), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n881), .B(new_n882), .C1(new_n201), .C2(new_n803), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(G50), .B2(new_n834), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n830), .A2(G87), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n822), .B2(new_n816), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT98), .Z(new_n888));
  INV_X1    g0688(.A(new_n824), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n450), .B1(new_n821), .B2(new_n506), .C1(new_n804), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G107), .B2(new_n834), .ZN(new_n891));
  AOI22_X1  g0691(.A1(G97), .A2(new_n843), .B1(new_n808), .B2(G283), .ZN(new_n892));
  INV_X1    g0692(.A(new_n813), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n891), .B(new_n892), .C1(new_n489), .C2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n885), .B1(new_n888), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n801), .B1(new_n895), .B2(KEYINPUT100), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(KEYINPUT100), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n797), .A2(new_n782), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n872), .B1(new_n898), .B2(new_n285), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n897), .B(new_n899), .C1(new_n783), .C2(new_n858), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n874), .A2(new_n900), .ZN(G384));
  NOR2_X1   g0701(.A1(new_n775), .A2(new_n211), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT16), .B1(new_n443), .B2(new_n453), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n420), .B1(new_n456), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n699), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n475), .A2(new_n476), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n479), .A3(new_n482), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(new_n469), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n473), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n907), .A3(new_n457), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n478), .A2(new_n473), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n478), .A2(new_n906), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n457), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n903), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n917), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n479), .A2(new_n482), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n468), .B1(new_n921), .B2(new_n908), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT38), .B(new_n920), .C1(new_n922), .C2(new_n907), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n377), .A2(new_n379), .A3(new_n701), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n363), .A2(new_n361), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n362), .B1(new_n358), .B2(G169), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n391), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n669), .A2(new_n925), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n380), .B2(new_n364), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n858), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n751), .A2(new_n759), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n751), .A2(KEYINPUT105), .A3(new_n759), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n752), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n932), .B1(new_n734), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT40), .B1(new_n924), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT104), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n457), .A2(new_n458), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT17), .B1(new_n466), .B2(new_n416), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n459), .A2(new_n467), .A3(KEYINPUT104), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n668), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n915), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n914), .A2(new_n915), .A3(new_n457), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n945), .A2(new_n946), .B1(new_n917), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n923), .B1(new_n949), .B2(KEYINPUT38), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n951), .B(new_n932), .C1(new_n734), .C2(new_n937), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n939), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n486), .B1(new_n734), .B2(new_n937), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n713), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT106), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(new_n953), .C2(new_n954), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n929), .A2(new_n931), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n852), .B(KEYINPUT103), .Z(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n868), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n924), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n482), .A2(new_n475), .A3(new_n699), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT39), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n945), .A2(new_n946), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n948), .A2(new_n917), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT38), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n910), .A2(new_n903), .A3(new_n918), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n364), .A2(new_n380), .A3(new_n702), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT39), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n485), .B1(new_n771), .B2(new_n772), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n672), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n978), .B(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n902), .B1(new_n960), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n960), .ZN(new_n983));
  INV_X1    g0783(.A(new_n600), .ZN(new_n984));
  OAI211_X1 g0784(.A(G116), .B(new_n227), .C1(new_n984), .C2(KEYINPUT35), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT102), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(KEYINPUT35), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(KEYINPUT102), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT36), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n793), .A2(G77), .A3(new_n447), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(G50), .B2(new_n202), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(G1), .A3(new_n280), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n983), .A2(new_n990), .A3(new_n993), .ZN(G367));
  NAND2_X1  g0794(.A1(new_n616), .A2(new_n701), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n610), .A2(new_n619), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT108), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n684), .A2(new_n701), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n723), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n649), .A2(new_n650), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n619), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n702), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n702), .A2(new_n675), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n565), .A3(new_n676), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n767), .B2(new_n1008), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT107), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(KEYINPUT43), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT109), .Z(new_n1015));
  AND3_X1   g0815(.A1(new_n1007), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1013), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n719), .A2(new_n999), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n726), .B(KEYINPUT41), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n723), .A2(new_n720), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n999), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT44), .Z(new_n1025));
  NOR2_X1   g0825(.A1(new_n999), .A2(new_n1023), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT45), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n719), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(new_n719), .A3(new_n1027), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n723), .B1(new_n718), .B2(new_n722), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n714), .B(new_n1031), .Z(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n773), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1022), .B1(new_n1033), .B2(new_n773), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1020), .B(new_n1021), .C1(new_n1034), .C2(new_n777), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n291), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n799), .B1(new_n725), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n791), .A2(new_n238), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n872), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(G283), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n821), .A2(new_n1040), .B1(new_n250), .B2(new_n803), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n809), .A2(new_n804), .B1(new_n893), .B2(new_n822), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n837), .C2(G303), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT46), .B1(new_n834), .B2(G116), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT110), .Z(new_n1045));
  NAND3_X1  g0845(.A1(new_n834), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n247), .B1(new_n817), .B2(G317), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n830), .A2(G97), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT111), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n803), .A2(new_n202), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n809), .B2(new_n437), .C1(new_n893), .C2(new_n877), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G50), .A2(new_n820), .B1(new_n824), .B2(G150), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n834), .A2(G58), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n830), .A2(G77), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n450), .B1(new_n817), .B2(G137), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT47), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n1039), .B1(new_n785), .B2(new_n1010), .C1(new_n1062), .C2(new_n801), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1035), .A2(new_n1063), .ZN(G387));
  AOI21_X1  g0864(.A(new_n727), .B1(new_n1032), .B2(new_n773), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n773), .B2(new_n1032), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n718), .A2(new_n785), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n791), .B1(new_n235), .B2(new_n538), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n729), .B2(new_n787), .ZN(new_n1069));
  OR3_X1    g0869(.A1(new_n309), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT50), .B1(new_n309), .B2(G50), .ZN(new_n1071));
  AOI21_X1  g0871(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n729), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1069), .A2(new_n1073), .B1(new_n250), .B2(new_n725), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n778), .B1(new_n1074), .B2(new_n799), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n437), .A2(new_n893), .B1(new_n809), .B2(new_n309), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n889), .A2(new_n317), .B1(new_n816), .B2(new_n310), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n247), .B1(new_n821), .B2(new_n202), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n834), .A2(G77), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n567), .A2(new_n843), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1079), .A2(new_n1048), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n837), .A2(G317), .B1(G303), .B2(new_n820), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G311), .A2(new_n808), .B1(new_n813), .B2(G322), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT113), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1040), .A2(new_n803), .B1(new_n833), .B2(new_n804), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(KEYINPUT49), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n247), .B1(new_n817), .B2(G326), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n506), .C2(new_n829), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT49), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1082), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1075), .B1(new_n1096), .B2(new_n797), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1032), .A2(new_n777), .B1(new_n1067), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1066), .A2(new_n1098), .ZN(G393));
  INV_X1    g0899(.A(new_n1030), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1100), .A2(new_n776), .A3(new_n1028), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n999), .A2(new_n784), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n798), .B1(new_n549), .B2(new_n218), .C1(new_n792), .C2(new_n245), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n778), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n809), .A2(new_n489), .B1(new_n506), .B2(new_n803), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n450), .B1(new_n821), .B2(new_n804), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G322), .C2(new_n817), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n250), .B2(new_n829), .C1(new_n1040), .C2(new_n833), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n824), .A2(G311), .B1(new_n813), .B2(G317), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n247), .B1(new_n821), .B2(new_n309), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n817), .B2(new_n878), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G77), .A2(new_n843), .B1(new_n808), .B2(G50), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n834), .A2(G68), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1113), .A2(new_n886), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n824), .A2(G159), .B1(new_n813), .B2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT51), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1108), .A2(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1104), .B1(new_n1119), .B2(new_n797), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1101), .B1(new_n1102), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1032), .A2(new_n773), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n1100), .B2(new_n1028), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1033), .A2(new_n1123), .A3(new_n726), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(G390));
  INV_X1    g0925(.A(G330), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n734), .B2(new_n937), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n485), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n979), .A2(new_n672), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n868), .A2(new_n962), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n961), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n761), .B2(new_n858), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1126), .B(new_n932), .C1(new_n734), .C2(new_n937), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n734), .A2(new_n760), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1135), .A2(new_n713), .A3(new_n858), .A4(new_n1131), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n861), .B1(new_n709), .B2(new_n1003), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n765), .A2(new_n768), .A3(new_n688), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n702), .B(new_n858), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n962), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1126), .B(new_n859), .C1(new_n734), .C2(new_n937), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1136), .B(new_n1141), .C1(new_n1142), .C2(new_n1131), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1129), .B1(new_n1134), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n975), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n973), .B2(new_n976), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1131), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n950), .A2(new_n1147), .A3(new_n974), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1133), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n974), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n468), .A2(new_n940), .B1(new_n475), .B2(new_n482), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n915), .B1(new_n1152), .B2(new_n944), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n970), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n903), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT39), .B1(new_n1155), .B2(new_n923), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n919), .A2(new_n923), .A3(KEYINPUT39), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1151), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n950), .A2(new_n1147), .A3(new_n974), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1136), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1144), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1149), .A2(new_n1160), .A3(new_n1144), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n726), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1149), .A2(new_n1160), .A3(new_n777), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n898), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n778), .B1(new_n1166), .B2(new_n295), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n450), .B1(new_n889), .B2(new_n506), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G294), .B2(new_n817), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G77), .A2(new_n843), .B1(new_n813), .B2(G283), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1169), .A2(new_n842), .A3(new_n882), .A4(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G97), .A2(new_n820), .B1(new_n808), .B2(G107), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT115), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n808), .A2(G137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n437), .B2(new_n803), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G128), .B2(new_n813), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n830), .A2(G50), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n450), .B1(new_n824), .B2(G132), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT54), .B(G143), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n820), .A2(new_n1180), .B1(new_n817), .B2(G125), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n834), .A2(G150), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT53), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1171), .A2(new_n1173), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1167), .B1(new_n1185), .B2(new_n797), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n783), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1165), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1164), .A2(new_n1190), .ZN(G378));
  AOI22_X1  g0991(.A1(G150), .A2(new_n843), .B1(new_n813), .B2(G125), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT116), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n834), .A2(new_n1180), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n808), .A2(G132), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G128), .A2(new_n824), .B1(new_n820), .B2(G137), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n817), .C2(G124), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n437), .B2(new_n829), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n247), .A2(G41), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n317), .B1(G33), .B2(G41), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1054), .B1(new_n549), .B2(new_n809), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G116), .B2(new_n813), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n824), .A2(G107), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n817), .A2(G283), .ZN(new_n1209));
  AND4_X1   g1009(.A1(new_n1080), .A2(new_n1208), .A3(new_n1209), .A4(new_n1203), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n567), .A2(new_n820), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n830), .A2(G58), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1207), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1205), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1214), .B2(new_n1213), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n797), .B1(new_n1202), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n778), .C1(G50), .C2(new_n1166), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n665), .A2(new_n333), .A3(new_n666), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n324), .A2(new_n699), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1220), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n665), .A2(new_n333), .A3(new_n666), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1221), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1218), .B1(new_n1230), .B2(new_n782), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n907), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n484), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT38), .B1(new_n1233), .B2(new_n920), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n938), .B1(new_n1234), .B2(new_n972), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n951), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1126), .B1(new_n950), .B2(new_n952), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1229), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1229), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n978), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n966), .B1(new_n1187), .B2(new_n975), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n971), .A2(new_n972), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n938), .A2(KEYINPUT40), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G330), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1230), .B1(new_n1244), .B2(new_n939), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1236), .A2(new_n1237), .A3(new_n1229), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1241), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1240), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1231), .B1(new_n1248), .B2(new_n777), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1241), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1245), .A2(new_n1246), .B1(new_n977), .B2(new_n967), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1129), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1163), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n726), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1163), .A2(new_n1253), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1249), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT117), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(KEYINPUT117), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(G375));
  NAND2_X1  g1065(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n777), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1166), .A2(G68), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n821), .A2(new_n310), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n450), .B(new_n1269), .C1(G128), .C2(new_n817), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n837), .A2(G137), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n834), .A2(G159), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1270), .A2(new_n1212), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G50), .A2(new_n843), .B1(new_n813), .B2(G132), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n809), .B2(new_n1179), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n450), .B1(new_n816), .B2(new_n489), .C1(new_n889), .C2(new_n1040), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G294), .B2(new_n813), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n834), .A2(G97), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1058), .A3(new_n1081), .A4(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(G107), .A2(new_n820), .B1(new_n808), .B2(G116), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT118), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1273), .A2(new_n1275), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n872), .B(new_n1268), .C1(new_n1282), .C2(new_n797), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1131), .B2(new_n783), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1267), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1144), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1022), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1134), .A2(new_n1129), .A3(new_n1143), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(G381));
  INV_X1    g1091(.A(G390), .ZN(new_n1292));
  INV_X1    g1092(.A(G384), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1066), .A2(new_n850), .A3(new_n1098), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1292), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(G387), .A3(G381), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1149), .A2(new_n1160), .A3(new_n1144), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1298), .A2(new_n1161), .A3(new_n727), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT119), .B1(new_n1299), .B2(new_n1189), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT119), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1164), .A2(new_n1301), .A3(new_n1190), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1297), .B(new_n1304), .C1(new_n1262), .C2(new_n1264), .ZN(G407));
  NOR2_X1   g1105(.A1(new_n694), .A2(G343), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G407), .B(G213), .C1(G375), .C2(new_n1307), .ZN(G409));
  INV_X1    g1108(.A(KEYINPUT126), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G378), .B(new_n1249), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1248), .A2(new_n1256), .A3(new_n1288), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1249), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1300), .A2(new_n1302), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1306), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT124), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(new_n1318), .A3(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1287), .A2(KEYINPUT60), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1320), .A2(new_n1289), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1134), .A2(new_n1129), .A3(new_n1143), .A4(KEYINPUT60), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n726), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G384), .B(new_n1286), .C1(new_n1321), .C2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1320), .B2(new_n1289), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1293), .B1(new_n1325), .B2(new_n1285), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1317), .A2(new_n1319), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1331), .B(new_n1328), .C1(new_n1316), .C2(new_n1327), .ZN(new_n1332));
  AOI211_X1 g1132(.A(new_n1306), .B(new_n1327), .C1(new_n1310), .C2(new_n1313), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1333), .B2(KEYINPUT62), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1330), .A2(new_n1332), .A3(new_n1334), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1336));
  INV_X1    g1136(.A(G2897), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1336), .A2(new_n1337), .A3(new_n1315), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT122), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT121), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1315), .B1(new_n1340), .B2(new_n1337), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1341), .B1(new_n1340), .B2(new_n1337), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1339), .B1(new_n1327), .B2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1336), .A2(KEYINPUT122), .A3(new_n1342), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1338), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1319), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1318), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1346), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT61), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1309), .B1(new_n1335), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n850), .B1(new_n1066), .B2(new_n1098), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1295), .A2(new_n1353), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1354), .A2(KEYINPUT123), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G387), .A2(new_n1292), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1035), .A2(G390), .A3(new_n1063), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1355), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  AND2_X1   g1158(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1354), .B(KEYINPUT123), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1358), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1330), .A2(new_n1332), .A3(new_n1334), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1362), .A2(KEYINPUT126), .A3(new_n1350), .A4(new_n1349), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1352), .A2(new_n1361), .A3(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1333), .A2(KEYINPUT63), .ZN(new_n1365));
  XOR2_X1   g1165(.A(new_n1365), .B(KEYINPUT120), .Z(new_n1366));
  AND2_X1   g1166(.A1(new_n1346), .A2(new_n1316), .ZN(new_n1367));
  NOR3_X1   g1167(.A1(new_n1367), .A2(new_n1361), .A3(KEYINPUT61), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1336), .A2(KEYINPUT63), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1366), .B(new_n1368), .C1(new_n1369), .C2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1364), .A2(new_n1371), .ZN(G405));
  NAND3_X1  g1172(.A1(new_n1261), .A2(new_n1263), .A3(new_n1304), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1373), .A2(new_n1310), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1375));
  XNOR2_X1  g1175(.A(new_n1374), .B(new_n1375), .ZN(new_n1376));
  XNOR2_X1  g1176(.A(new_n1376), .B(new_n1361), .ZN(G402));
endmodule


