

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U327 ( .A(n468), .B(KEYINPUT96), .ZN(n469) );
  XOR2_X1 U328 ( .A(G92GAT), .B(G64GAT), .Z(n350) );
  XNOR2_X1 U329 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U330 ( .A(G190GAT), .B(KEYINPUT78), .Z(n295) );
  XOR2_X1 U331 ( .A(n317), .B(n316), .Z(n543) );
  XNOR2_X1 U332 ( .A(n381), .B(KEYINPUT109), .ZN(n382) );
  XNOR2_X1 U333 ( .A(n383), .B(n382), .ZN(n399) );
  XNOR2_X1 U334 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U335 ( .A(n409), .B(KEYINPUT48), .ZN(n410) );
  XNOR2_X1 U336 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U337 ( .A(n350), .B(n295), .ZN(n339) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G85GAT), .Z(n362) );
  XNOR2_X1 U339 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n478) );
  XNOR2_X1 U340 ( .A(n340), .B(n339), .ZN(n344) );
  XNOR2_X1 U341 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U342 ( .A(n479), .B(n478), .ZN(n517) );
  XNOR2_X1 U343 ( .A(n364), .B(n363), .ZN(n579) );
  INV_X1 U344 ( .A(G190GAT), .ZN(n456) );
  INV_X1 U345 ( .A(G43GAT), .ZN(n483) );
  XNOR2_X1 U346 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U347 ( .A(n483), .B(KEYINPUT40), .ZN(n484) );
  XNOR2_X1 U348 ( .A(n485), .B(n484), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(n362), .B(G218GAT), .Z(n297) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G134GAT), .Z(n440) );
  XNOR2_X1 U351 ( .A(n440), .B(G162GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n299) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G92GAT), .ZN(n298) );
  XOR2_X1 U355 ( .A(n299), .B(n298), .Z(n301) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XOR2_X1 U357 ( .A(KEYINPUT75), .B(KEYINPUT73), .Z(n305) );
  XNOR2_X1 U358 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U360 ( .A(n307), .B(n306), .Z(n317) );
  XOR2_X1 U361 ( .A(G29GAT), .B(KEYINPUT7), .Z(n309) );
  XNOR2_X1 U362 ( .A(G50GAT), .B(G36GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U364 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n310) );
  XOR2_X1 U365 ( .A(n311), .B(n310), .Z(n379) );
  INV_X1 U366 ( .A(n379), .ZN(n315) );
  XOR2_X1 U367 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n313) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U370 ( .A(n315), .B(n314), .Z(n316) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G22GAT), .Z(n370) );
  XOR2_X1 U372 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n319) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(KEYINPUT88), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U375 ( .A(n370), .B(n320), .Z(n322) );
  NAND2_X1 U376 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n335) );
  XOR2_X1 U378 ( .A(G211GAT), .B(KEYINPUT24), .Z(n324) );
  XNOR2_X1 U379 ( .A(G78GAT), .B(KEYINPUT23), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n327) );
  XOR2_X1 U381 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n326) );
  XNOR2_X1 U382 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n336) );
  XOR2_X1 U384 ( .A(n327), .B(n336), .Z(n333) );
  XOR2_X1 U385 ( .A(KEYINPUT2), .B(G162GAT), .Z(n329) );
  XNOR2_X1 U386 ( .A(KEYINPUT90), .B(G155GAT), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U388 ( .A(KEYINPUT3), .B(n330), .Z(n424) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(G204GAT), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n331), .B(G148GAT), .ZN(n358) );
  XNOR2_X1 U391 ( .A(n424), .B(n358), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U393 ( .A(n335), .B(n334), .Z(n466) );
  XOR2_X1 U394 ( .A(KEYINPUT94), .B(n336), .Z(n338) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U397 ( .A(G204GAT), .B(G183GAT), .Z(n342) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G36GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U401 ( .A(G176GAT), .B(KEYINPUT19), .Z(n346) );
  XNOR2_X1 U402 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n449) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(G211GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n347), .B(KEYINPUT79), .ZN(n395) );
  XNOR2_X1 U406 ( .A(n449), .B(n395), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n521) );
  XNOR2_X1 U408 ( .A(G176GAT), .B(G120GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U410 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n353) );
  XNOR2_X1 U411 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U413 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U414 ( .A(KEYINPUT13), .B(G57GAT), .Z(n357) );
  XNOR2_X1 U415 ( .A(G71GAT), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n394) );
  XNOR2_X1 U417 ( .A(n358), .B(n394), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n364) );
  NAND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT41), .B(n579), .Z(n566) );
  XOR2_X1 U421 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n366) );
  XNOR2_X1 U422 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n378) );
  XOR2_X1 U424 ( .A(G8GAT), .B(G1GAT), .Z(n368) );
  XNOR2_X1 U425 ( .A(G197GAT), .B(G15GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U427 ( .A(n370), .B(n369), .Z(n372) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U430 ( .A(n373), .B(KEYINPUT29), .Z(n376) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G43GAT), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n374), .B(G113GAT), .ZN(n441) );
  XNOR2_X1 U433 ( .A(n441), .B(KEYINPUT30), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U436 ( .A(n380), .B(n379), .Z(n549) );
  INV_X1 U437 ( .A(n549), .ZN(n575) );
  NOR2_X1 U438 ( .A1(n566), .A2(n575), .ZN(n383) );
  XNOR2_X1 U439 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n381) );
  XOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n389) );
  XNOR2_X1 U441 ( .A(G15GAT), .B(G183GAT), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n384), .B(G127GAT), .ZN(n450) );
  XOR2_X1 U443 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n386) );
  XNOR2_X1 U444 ( .A(G1GAT), .B(G64GAT), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n450), .B(n387), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U448 ( .A(G155GAT), .B(G22GAT), .Z(n391) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U451 ( .A(n393), .B(n392), .Z(n397) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U453 ( .A(n397), .B(n396), .Z(n556) );
  XOR2_X1 U454 ( .A(KEYINPUT108), .B(n556), .Z(n570) );
  INV_X1 U455 ( .A(n543), .ZN(n558) );
  AND2_X1 U456 ( .A1(n570), .A2(n543), .ZN(n398) );
  AND2_X1 U457 ( .A1(n399), .A2(n398), .ZN(n401) );
  XNOR2_X1 U458 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n408) );
  INV_X1 U460 ( .A(n579), .ZN(n480) );
  INV_X1 U461 ( .A(n556), .ZN(n584) );
  XOR2_X1 U462 ( .A(n543), .B(KEYINPUT101), .Z(n402) );
  XNOR2_X1 U463 ( .A(n402), .B(KEYINPUT36), .ZN(n587) );
  NOR2_X1 U464 ( .A1(n584), .A2(n587), .ZN(n404) );
  XNOR2_X1 U465 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U467 ( .A(KEYINPUT71), .B(n575), .Z(n561) );
  NAND2_X1 U468 ( .A1(n405), .A2(n561), .ZN(n406) );
  NOR2_X1 U469 ( .A1(n480), .A2(n406), .ZN(n407) );
  NOR2_X1 U470 ( .A1(n408), .A2(n407), .ZN(n411) );
  INV_X1 U471 ( .A(KEYINPUT113), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n530) );
  NOR2_X1 U473 ( .A1(n521), .A2(n530), .ZN(n413) );
  XNOR2_X1 U474 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n435) );
  XOR2_X1 U476 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n415) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n417) );
  XNOR2_X1 U480 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U482 ( .A(n419), .B(n418), .Z(n426) );
  XNOR2_X1 U483 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n420), .B(KEYINPUT82), .ZN(n444) );
  XOR2_X1 U485 ( .A(n444), .B(KEYINPUT92), .Z(n422) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n434) );
  XOR2_X1 U490 ( .A(G148GAT), .B(G127GAT), .Z(n428) );
  XNOR2_X1 U491 ( .A(G113GAT), .B(G141GAT), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U493 ( .A(G85GAT), .B(KEYINPUT76), .Z(n430) );
  XNOR2_X1 U494 ( .A(G29GAT), .B(G134GAT), .ZN(n429) );
  XNOR2_X1 U495 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U496 ( .A(n432), .B(n431), .Z(n433) );
  XOR2_X1 U497 ( .A(n434), .B(n433), .Z(n460) );
  INV_X1 U498 ( .A(n460), .ZN(n519) );
  NAND2_X1 U499 ( .A1(n435), .A2(n519), .ZN(n436) );
  XOR2_X1 U500 ( .A(KEYINPUT64), .B(n436), .Z(n574) );
  NAND2_X1 U501 ( .A1(n466), .A2(n574), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n437), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U503 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n439) );
  XNOR2_X1 U504 ( .A(G71GAT), .B(KEYINPUT65), .ZN(n438) );
  XNOR2_X1 U505 ( .A(n439), .B(n438), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT85), .B(n440), .Z(n443) );
  XNOR2_X1 U507 ( .A(n441), .B(G99GAT), .ZN(n442) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n448) );
  XOR2_X1 U509 ( .A(n444), .B(KEYINPUT20), .Z(n446) );
  NAND2_X1 U510 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U512 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U514 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X2 U515 ( .A(n454), .B(n453), .Z(n523) );
  INV_X1 U516 ( .A(n523), .ZN(n531) );
  NAND2_X1 U517 ( .A1(n455), .A2(n531), .ZN(n569) );
  NOR2_X1 U518 ( .A1(n543), .A2(n569), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U521 ( .A(n523), .B(KEYINPUT86), .Z(n463) );
  XOR2_X1 U522 ( .A(n466), .B(KEYINPUT28), .Z(n497) );
  XOR2_X1 U523 ( .A(n521), .B(KEYINPUT27), .Z(n465) );
  NAND2_X1 U524 ( .A1(n460), .A2(n465), .ZN(n529) );
  NOR2_X1 U525 ( .A1(n497), .A2(n529), .ZN(n461) );
  XNOR2_X1 U526 ( .A(KEYINPUT95), .B(n461), .ZN(n462) );
  NOR2_X1 U527 ( .A1(n463), .A2(n462), .ZN(n476) );
  NOR2_X1 U528 ( .A1(n531), .A2(n466), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n464), .B(KEYINPUT26), .ZN(n573) );
  NAND2_X1 U530 ( .A1(n573), .A2(n465), .ZN(n472) );
  OR2_X1 U531 ( .A1(n523), .A2(n521), .ZN(n467) );
  NAND2_X1 U532 ( .A1(n467), .A2(n466), .ZN(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n468) );
  NAND2_X1 U534 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n473), .A2(n519), .ZN(n474) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(n474), .Z(n475) );
  NOR2_X1 U537 ( .A1(n476), .A2(n475), .ZN(n489) );
  NOR2_X1 U538 ( .A1(n587), .A2(n489), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n584), .A2(n477), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n561), .A2(n480), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n517), .A2(n490), .ZN(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT103), .B(n481), .Z(n482) );
  XNOR2_X1 U543 ( .A(KEYINPUT38), .B(n482), .ZN(n505) );
  NOR2_X1 U544 ( .A1(n523), .A2(n505), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n487) );
  NAND2_X1 U546 ( .A1(n556), .A2(n543), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n507) );
  NAND2_X1 U549 ( .A1(n490), .A2(n507), .ZN(n498) );
  NOR2_X1 U550 ( .A1(n519), .A2(n498), .ZN(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(n491), .Z(n492) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n521), .A2(n498), .ZN(n493) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n523), .A2(n498), .ZN(n495) );
  XNOR2_X1 U556 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  INV_X1 U559 ( .A(n497), .ZN(n533) );
  NOR2_X1 U560 ( .A1(n533), .A2(n498), .ZN(n499) );
  XOR2_X1 U561 ( .A(KEYINPUT100), .B(n499), .Z(n500) );
  XNOR2_X1 U562 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  NOR2_X1 U563 ( .A1(n505), .A2(n519), .ZN(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n521), .A2(n505), .ZN(n504) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U569 ( .A1(n505), .A2(n533), .ZN(n506) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  NOR2_X1 U571 ( .A1(n549), .A2(n566), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n518), .A2(n507), .ZN(n514) );
  NOR2_X1 U573 ( .A1(n519), .A2(n514), .ZN(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n521), .A2(n514), .ZN(n511) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n511), .Z(n512) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n523), .A2(n514), .ZN(n513) );
  XOR2_X1 U581 ( .A(G71GAT), .B(n513), .Z(G1334GAT) );
  NOR2_X1 U582 ( .A1(n533), .A2(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U586 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n525), .ZN(n524) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n533), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n547), .A2(n531), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT114), .B(n532), .Z(n534) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n561), .A2(n542), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  NOR2_X1 U603 ( .A1(n566), .A2(n542), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n570), .A2(n542), .ZN(n540) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n540), .Z(n541) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  NAND2_X1 U614 ( .A1(n573), .A2(n547), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(n548), .Z(n559) );
  NAND2_X1 U616 ( .A1(n549), .A2(n559), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .Z(n553) );
  INV_X1 U619 ( .A(n566), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n551), .A2(n559), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n556), .A2(n559), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n569), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n565) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n566), .ZN(n567) );
  XOR2_X1 U635 ( .A(n568), .B(n567), .Z(G1349GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n575), .A2(n586), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n586), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

