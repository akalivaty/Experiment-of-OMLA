//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT22), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT75), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n210), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT76), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(KEYINPUT75), .B2(new_n211), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n212), .B1(new_n209), .B2(new_n208), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI221_X1 g024(.A(new_n220), .B1(KEYINPUT68), .B2(KEYINPUT28), .C1(new_n221), .C2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(G169gat), .ZN(new_n230));
  INV_X1    g029(.A(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT26), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(KEYINPUT26), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n229), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n239), .A2(G169gat), .A3(G176gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n234), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n229), .ZN(new_n244));
  AND2_X1   g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT24), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(KEYINPUT67), .B(new_n234), .C1(new_n232), .C2(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n239), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n242), .A2(new_n247), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT25), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G176gat), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n239), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT65), .B(G169gat), .Z(new_n256));
  AOI21_X1  g055(.A(KEYINPUT25), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n241), .B1(new_n239), .B2(new_n232), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(KEYINPUT64), .A3(KEYINPUT24), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n246), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n257), .A2(new_n258), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n237), .A2(new_n251), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n219), .B(new_n265), .C1(new_n267), .C2(new_n264), .ZN(new_n268));
  INV_X1    g067(.A(new_n219), .ZN(new_n269));
  INV_X1    g068(.A(new_n265), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n264), .B1(new_n263), .B2(new_n266), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274));
  INV_X1    g073(.A(G64gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n273), .B2(new_n278), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n279), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G78gat), .B(G106gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT84), .B(G22gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT2), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G141gat), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G148gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n288), .B(new_n290), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G155gat), .B(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(G141gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT77), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n296), .A3(new_n290), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n286), .A3(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n266), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n214), .A2(new_n218), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G228gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n308), .B(KEYINPUT85), .ZN(new_n312));
  INV_X1    g111(.A(new_n211), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT29), .B1(new_n210), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n313), .B2(new_n210), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n286), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n303), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n307), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n285), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n285), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n307), .A2(new_n317), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n320), .B(new_n310), .C1(new_n321), .C2(new_n312), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT31), .B(G50gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n319), .B2(new_n322), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G113gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G120gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G127gat), .B(G134gat), .Z(new_n337));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n337), .B1(KEYINPUT1), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n263), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n339), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n237), .A2(new_n262), .A3(new_n251), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT34), .ZN(new_n345));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT34), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n344), .A2(KEYINPUT71), .A3(new_n345), .A4(new_n346), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n346), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n341), .A2(new_n354), .A3(new_n343), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT33), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G15gat), .B(G43gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G71gat), .ZN(new_n360));
  INV_X1    g159(.A(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(KEYINPUT33), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(KEYINPUT32), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n353), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n353), .A2(new_n366), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(KEYINPUT87), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n282), .B(new_n326), .C1(new_n370), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n302), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n296), .B1(new_n301), .B2(new_n290), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n342), .A3(new_n305), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n298), .A4(new_n302), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n298), .A2(new_n336), .A3(new_n302), .A4(new_n339), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n303), .A2(new_n342), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n380), .ZN(new_n387));
  INV_X1    g186(.A(new_n379), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT79), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n390));
  AOI211_X1 g189(.A(new_n390), .B(new_n379), .C1(new_n386), .C2(new_n380), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n384), .B(new_n385), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n380), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n381), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n385), .A2(new_n388), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n394), .A2(new_n377), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G57gat), .ZN(new_n401));
  INV_X1    g200(.A(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AND4_X1   g203(.A1(KEYINPUT82), .A2(new_n398), .A3(KEYINPUT6), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n392), .B2(new_n397), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT82), .B1(new_n406), .B2(KEYINPUT6), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n398), .A2(new_n404), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n403), .A3(new_n397), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n413), .A2(KEYINPUT35), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n373), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT70), .ZN(new_n416));
  INV_X1    g215(.A(new_n365), .ZN(new_n417));
  INV_X1    g216(.A(new_n362), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n355), .B2(new_n357), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n363), .A2(KEYINPUT70), .A3(new_n365), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n422), .A2(new_n423), .A3(new_n353), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n422), .B2(new_n353), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n426), .A2(KEYINPUT88), .A3(new_n326), .A4(new_n367), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT81), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n409), .A2(new_n429), .A3(new_n411), .A4(new_n410), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n408), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n273), .A2(new_n278), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n281), .B(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT83), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n417), .A2(new_n419), .A3(new_n416), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT70), .B1(new_n363), .B2(new_n365), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n353), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n353), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n326), .A3(new_n367), .A4(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n408), .A2(new_n428), .A3(new_n430), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n282), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n427), .A2(new_n434), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n415), .B1(new_n446), .B2(KEYINPUT35), .ZN(new_n447));
  INV_X1    g246(.A(new_n326), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n443), .A2(new_n444), .A3(new_n282), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n443), .B2(new_n282), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT36), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n369), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT73), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n438), .A2(KEYINPUT36), .A3(new_n367), .A4(new_n439), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n369), .A2(new_n456), .A3(new_n452), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT37), .B1(new_n273), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n268), .A2(new_n272), .A3(KEYINPUT86), .A4(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n278), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n432), .B1(new_n463), .B2(KEYINPUT38), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT38), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n460), .A2(new_n465), .A3(new_n278), .A4(new_n462), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n464), .A2(new_n408), .A3(new_n412), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n394), .A2(new_n377), .A3(new_n395), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n388), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n469), .B(KEYINPUT39), .C1(new_n388), .C2(new_n387), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n470), .B(new_n403), .C1(KEYINPUT39), .C2(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n433), .A2(new_n473), .A3(new_n409), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n467), .A2(new_n475), .A3(new_n326), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n451), .A2(new_n458), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n447), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G231gat), .ZN(new_n479));
  INV_X1    g278(.A(G233gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n275), .A2(G57gat), .ZN(new_n482));
  INV_X1    g281(.A(G57gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G64gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT94), .ZN(new_n486));
  NAND2_X1  g285(.A1(G71gat), .A2(G78gat), .ZN(new_n487));
  OR2_X1    g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT9), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n482), .A2(new_n484), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT9), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n487), .A3(new_n488), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n491), .A2(new_n496), .A3(KEYINPUT95), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT95), .B1(new_n491), .B2(new_n496), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G127gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n503), .A2(G127gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n481), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  INV_X1    g307(.A(new_n481), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n514), .A2(KEYINPUT91), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n514), .B2(KEYINPUT91), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n514), .A2(KEYINPUT16), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n514), .A2(new_n515), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n520), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n498), .A2(KEYINPUT21), .A3(new_n500), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT96), .B(G155gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n526), .A2(new_n527), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(new_n528), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n529), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(new_n510), .A3(new_n507), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n536));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n534), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n544), .A2(G29gat), .A3(G36gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G29gat), .A2(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT14), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n546), .B1(KEYINPUT14), .B2(new_n548), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(new_n545), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G43gat), .B(G50gat), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n550), .B2(KEYINPUT15), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n556), .B1(new_n551), .B2(new_n554), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT89), .B1(new_n563), .B2(new_n560), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n566), .B1(new_n558), .B2(new_n561), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n570), .A2(KEYINPUT97), .B1(KEYINPUT8), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n402), .A2(new_n277), .ZN(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT7), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n570), .A2(KEYINPUT97), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n567), .A2(new_n569), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n576), .B(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT98), .ZN(new_n586));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n580), .A2(new_n588), .A3(new_n582), .A4(new_n584), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n586), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n543), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n589), .ZN(new_n593));
  INV_X1    g392(.A(new_n587), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(KEYINPUT99), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n592), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n543), .B(new_n600), .C1(new_n590), .C2(new_n591), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT100), .B1(new_n542), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n542), .A2(new_n604), .A3(KEYINPUT100), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n478), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n568), .B1(new_n565), .B2(new_n566), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n526), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n523), .A2(new_n525), .A3(new_n565), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n608), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n565), .B1(new_n523), .B2(new_n525), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n611), .A4(new_n613), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n615), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT11), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n230), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n579), .B1(new_n497), .B2(new_n499), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n491), .A2(new_n496), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n581), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n498), .A2(new_n500), .A3(new_n581), .A4(KEYINPUT10), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n231), .ZN(new_n643));
  INV_X1    g442(.A(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n640), .B1(new_n632), .B2(new_n636), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT101), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n645), .B(KEYINPUT102), .Z(new_n652));
  INV_X1    g451(.A(new_n641), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n648), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n631), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n607), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n431), .A2(KEYINPUT103), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n431), .A2(KEYINPUT103), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n515), .ZN(G1324gat));
  INV_X1    g462(.A(new_n657), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n433), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT16), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n520), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n666), .A2(new_n668), .B1(G8gat), .B2(new_n665), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n670), .ZN(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n657), .A2(new_n674), .A3(new_n458), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n370), .A2(new_n372), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n664), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n674), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n657), .A2(new_n326), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  AND2_X1   g480(.A1(new_n602), .A2(new_n603), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n451), .A2(KEYINPUT105), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n458), .A2(new_n476), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n685), .B(new_n448), .C1(new_n449), .C2(new_n450), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n687), .B2(new_n447), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n655), .B(KEYINPUT104), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n542), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n682), .C1(new_n447), .C2(new_n477), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n690), .A2(new_n630), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n661), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n478), .A2(new_n604), .ZN(new_n697));
  INV_X1    g496(.A(new_n542), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n656), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(G29gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n696), .B1(new_n700), .B2(new_n660), .ZN(new_n701));
  NOR4_X1   g500(.A1(new_n699), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n661), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n695), .B1(new_n701), .B2(new_n702), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n699), .A2(G36gat), .A3(new_n282), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n706), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n694), .A2(new_n282), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT107), .Z(new_n710));
  INV_X1    g509(.A(G36gat), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n707), .B(new_n708), .C1(new_n710), .C2(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(G43gat), .B1(new_n694), .B2(new_n458), .ZN(new_n713));
  INV_X1    g512(.A(new_n676), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n699), .A2(G43gat), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT108), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g516(.A(G50gat), .B1(new_n694), .B2(new_n326), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n326), .A2(G50gat), .ZN(new_n719));
  OAI221_X1 g518(.A(new_n718), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n699), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n723));
  INV_X1    g522(.A(new_n415), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n606), .A2(new_n605), .A3(new_n630), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n727), .A2(new_n691), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n660), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n433), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  AOI21_X1  g534(.A(G71gat), .B1(new_n729), .B2(new_n676), .ZN(new_n736));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n458), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n729), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g539(.A1(new_n729), .A2(new_n448), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G78gat), .ZN(G1335gat));
  INV_X1    g541(.A(new_n655), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n542), .A2(new_n630), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n604), .B1(new_n725), .B2(new_n726), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n693), .B(new_n744), .C1(new_n745), .C2(KEYINPUT44), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n661), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n727), .A2(new_n631), .A3(new_n698), .A4(new_n682), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT111), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n655), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n660), .A2(new_n402), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(G1336gat));
  OAI211_X1 g555(.A(KEYINPUT112), .B(G92gat), .C1(new_n748), .C2(new_n282), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n690), .A2(new_n747), .A3(new_n693), .A4(new_n744), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n746), .A2(KEYINPUT110), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n282), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(new_n277), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n752), .A2(new_n277), .A3(new_n433), .A4(new_n691), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n757), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n746), .B2(new_n282), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n748), .B2(new_n458), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n676), .A2(new_n361), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n754), .B2(new_n771), .ZN(G1338gat));
  INV_X1    g571(.A(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n691), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n326), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n752), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n752), .A2(KEYINPUT114), .A3(new_n773), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT113), .B(G106gat), .Z(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n748), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n448), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT53), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n781), .B1(new_n746), .B2(new_n326), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n776), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n637), .A2(G230gat), .A3(G233gat), .A4(new_n638), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n641), .A2(KEYINPUT54), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n641), .A2(new_n795), .A3(KEYINPUT54), .A4(new_n791), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n793), .A2(new_n645), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT55), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n646), .B1(new_n792), .B2(KEYINPUT115), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n794), .A4(new_n796), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n630), .A2(new_n802), .A3(new_n651), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n612), .A2(new_n614), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT116), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n618), .A2(new_n619), .A3(new_n617), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n612), .A2(new_n807), .A3(new_n614), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n627), .A2(new_n622), .B1(new_n809), .B2(new_n626), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n655), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n682), .B1(new_n803), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n650), .B1(new_n798), .B2(new_n801), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n602), .A2(new_n810), .A3(new_n603), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n790), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n682), .A2(new_n810), .A3(new_n813), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n813), .A2(new_n630), .B1(new_n655), .B2(new_n810), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n818), .B(KEYINPUT117), .C1(new_n819), .C2(new_n682), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n698), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n728), .A2(new_n743), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n661), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n427), .A2(new_n442), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n823), .A2(new_n282), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n329), .A3(new_n630), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n660), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n631), .A3(new_n373), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n329), .B2(new_n829), .ZN(G1340gat));
  NOR2_X1   g629(.A1(new_n828), .A2(new_n373), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n691), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n655), .A2(new_n327), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT118), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n832), .A2(G120gat), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT119), .ZN(G1341gat));
  AOI21_X1  g635(.A(G127gat), .B1(new_n825), .B2(new_n542), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n542), .A2(G127gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n831), .B2(new_n838), .ZN(G1342gat));
  NAND2_X1  g638(.A1(new_n831), .A2(new_n682), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G134gat), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n282), .A3(new_n824), .A4(new_n682), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT56), .B1(new_n842), .B2(G134gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT120), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n841), .A2(new_n843), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1343gat));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n827), .A2(new_n850), .A3(new_n448), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n818), .B1(new_n819), .B2(new_n682), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n728), .A2(new_n743), .B1(new_n852), .B2(new_n698), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT57), .B1(new_n853), .B2(new_n326), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n660), .A2(new_n282), .A3(new_n458), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n851), .A2(new_n630), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G141gat), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT58), .B1(new_n858), .B2(KEYINPUT122), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n828), .A2(KEYINPUT121), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n458), .A2(new_n448), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n282), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n823), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n631), .A2(G141gat), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n860), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n858), .B(new_n866), .C1(KEYINPUT122), .C2(KEYINPUT58), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1344gat));
  AND3_X1   g669(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n291), .A3(new_n655), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n851), .A2(new_n854), .A3(new_n856), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n743), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n291), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n827), .A2(KEYINPUT57), .A3(new_n448), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n850), .B1(new_n853), .B2(new_n326), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n655), .A3(new_n856), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(G148gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n872), .B1(new_n876), .B2(new_n881), .ZN(G1345gat));
  INV_X1    g681(.A(G155gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n874), .A2(new_n883), .A3(new_n698), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n871), .A2(new_n542), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n883), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n887), .A3(new_n682), .ZN(new_n888));
  OAI21_X1  g687(.A(G162gat), .B1(new_n874), .B2(new_n604), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1347gat));
  AOI21_X1  g689(.A(new_n660), .B1(new_n821), .B2(new_n822), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(new_n433), .A3(new_n824), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n630), .A3(new_n256), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n660), .A2(new_n282), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n676), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT123), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n827), .A2(new_n326), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n631), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT124), .Z(G1348gat));
  AOI21_X1  g699(.A(G176gat), .B1(new_n892), .B2(new_n655), .ZN(new_n901));
  INV_X1    g700(.A(new_n897), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n691), .A2(new_n252), .A3(new_n254), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(G1349gat));
  OAI211_X1 g703(.A(new_n892), .B(new_n542), .C1(new_n222), .C2(new_n221), .ZN(new_n905));
  OAI21_X1  g704(.A(G183gat), .B1(new_n897), .B2(new_n698), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n897), .B2(new_n604), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT61), .B1(new_n909), .B2(KEYINPUT126), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n220), .A3(new_n682), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n879), .A2(new_n458), .A3(new_n894), .ZN(new_n918));
  OAI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n631), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n891), .A2(new_n433), .A3(new_n861), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n631), .A2(G197gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  NOR3_X1   g721(.A1(new_n920), .A2(G204gat), .A3(new_n743), .ZN(new_n923));
  XNOR2_X1  g722(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G204gat), .B1(new_n918), .B2(new_n774), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G1353gat));
  INV_X1    g728(.A(new_n920), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n206), .A3(new_n542), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n879), .A2(new_n458), .A3(new_n542), .A4(new_n894), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n207), .A3(new_n604), .ZN(new_n936));
  AOI21_X1  g735(.A(G218gat), .B1(new_n930), .B2(new_n682), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


