//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n204));
  OR3_X1    g003(.A1(new_n203), .A2(new_n204), .A3(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n205), .B(new_n207), .C1(new_n209), .C2(G8gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215));
  INV_X1    g014(.A(G71gat), .ZN(new_n216));
  INV_X1    g015(.A(G78gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(KEYINPUT95), .ZN(new_n221));
  INV_X1    g020(.A(G57gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G64gat), .ZN(new_n223));
  INV_X1    g022(.A(G64gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G57gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n221), .B(new_n226), .Z(new_n227));
  OAI21_X1  g026(.A(new_n214), .B1(new_n215), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n229));
  NAND2_X1  g028(.A1(G231gat), .A2(G233gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n228), .B(new_n231), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n215), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT96), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n235), .A2(KEYINPUT97), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(KEYINPUT97), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G155gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT20), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G183gat), .B(G211gat), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n240), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n244), .A3(new_n237), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n241), .B2(new_n245), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n233), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n242), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n232), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G218gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n255), .A2(KEYINPUT15), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(G29gat), .B2(G36gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(G29gat), .A2(G36gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT14), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n257), .B(new_n260), .C1(KEYINPUT15), .C2(new_n255), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(KEYINPUT90), .ZN(new_n262));
  NAND2_X1  g061(.A1(G29gat), .A2(G36gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n256), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT17), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(KEYINPUT17), .A3(new_n266), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT102), .B(G92gat), .Z(new_n271));
  INV_X1    g070(.A(G85gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G99gat), .A2(G106gat), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n271), .A2(new_n272), .B1(KEYINPUT8), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT101), .B(KEYINPUT7), .ZN(new_n275));
  NAND3_X1  g074(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n276), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G99gat), .B(G106gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n274), .A2(new_n277), .A3(new_n280), .A4(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n270), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n284), .ZN(new_n287));
  AND2_X1   g086(.A1(G232gat), .A2(G233gat), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(new_n267), .B1(KEYINPUT41), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n286), .B1(new_n285), .B2(new_n289), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n254), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(G218gat), .A3(new_n290), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT99), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n288), .A2(KEYINPUT41), .ZN(new_n298));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(new_n300), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT103), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n253), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n248), .A2(new_n252), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT103), .B1(new_n308), .B2(new_n304), .ZN(new_n309));
  XNOR2_X1  g108(.A(G120gat), .B(G148gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  XOR2_X1   g111(.A(new_n312), .B(KEYINPUT104), .Z(new_n313));
  NAND2_X1  g112(.A1(new_n284), .A2(new_n227), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n221), .B(new_n226), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n282), .A2(new_n316), .A3(new_n283), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G230gat), .A2(G233gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT105), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT105), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n325), .A3(new_n322), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n314), .B2(new_n317), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n313), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n330), .A3(new_n312), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n307), .A2(new_n309), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G127gat), .ZN(new_n337));
  INV_X1    g136(.A(G127gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G134gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n337), .A2(new_n339), .B1(new_n340), .B2(G134gat), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT72), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n336), .A2(KEYINPUT71), .ZN(new_n346));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G113gat), .B(G120gat), .Z(new_n349));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n353), .A3(new_n347), .ZN(new_n354));
  INV_X1    g153(.A(G141gat), .ZN(new_n355));
  INV_X1    g154(.A(G148gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n361));
  INV_X1    g160(.A(G155gat), .ZN(new_n362));
  INV_X1    g161(.A(G162gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n359), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(KEYINPUT2), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT79), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(G155gat), .B2(G162gat), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n369), .A2(new_n371), .A3(new_n360), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n366), .A2(new_n357), .A3(new_n358), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n365), .A2(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n354), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n352), .A2(new_n374), .A3(new_n377), .A4(new_n354), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n335), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT5), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n373), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n360), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(new_n368), .A3(new_n357), .A4(new_n358), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n354), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n344), .B1(new_n347), .B2(new_n346), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n393), .A2(KEYINPUT72), .B1(new_n350), .B2(new_n349), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n394), .B2(new_n348), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n382), .B(new_n383), .C1(new_n391), .C2(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n379), .A2(new_n381), .A3(new_n396), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT82), .B(new_n374), .C1(new_n352), .C2(new_n354), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n352), .A2(new_n354), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n387), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n376), .B(new_n378), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n383), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n382), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n391), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n376), .A2(new_n335), .A3(new_n378), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n397), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  AOI21_X1  g213(.A(KEYINPUT6), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n401), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n376), .A2(new_n378), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n403), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT5), .A3(new_n409), .ZN(new_n419));
  INV_X1    g218(.A(new_n397), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n410), .A2(KEYINPUT86), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n414), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n410), .B2(KEYINPUT86), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n422), .B(new_n397), .C1(new_n404), .C2(new_n409), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n415), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n432), .B(new_n414), .C1(new_n419), .C2(new_n420), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G197gat), .B(G204gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT22), .ZN(new_n436));
  INV_X1    g235(.A(G211gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n254), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G211gat), .B(G218gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n435), .A3(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT26), .ZN(new_n449));
  NAND2_X1  g248(.A1(G183gat), .A2(G190gat), .ZN(new_n450));
  INV_X1    g249(.A(G169gat), .ZN(new_n451));
  INV_X1    g250(.A(G176gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT26), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT69), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G190gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT27), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G183gat), .ZN(new_n461));
  INV_X1    g260(.A(G183gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT27), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n457), .A2(new_n459), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT28), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT68), .B(G183gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT27), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT69), .B(G190gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT28), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT70), .B1(new_n462), .B2(KEYINPUT27), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT70), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n460), .A3(G183gat), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n456), .B(new_n465), .C1(new_n468), .C2(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT24), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n450), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT65), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n286), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT23), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(G176gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n446), .A2(KEYINPUT23), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n489), .A2(new_n491), .B1(new_n453), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n477), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT23), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n490), .B1(G169gat), .B2(G176gat), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT25), .B(new_n495), .C1(new_n496), .C2(new_n448), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n478), .A2(new_n462), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n466), .A2(new_n469), .B1(G190gat), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT24), .B1(new_n450), .B2(KEYINPUT67), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(KEYINPUT67), .B2(new_n450), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n475), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n503), .A2(new_n504), .B1(G226gat), .B2(G233gat), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n485), .B(new_n482), .C1(new_n483), .C2(KEYINPUT65), .ZN(new_n506));
  INV_X1    g305(.A(new_n484), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT66), .B(G169gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n491), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n509), .A2(new_n510), .B1(new_n496), .B2(new_n448), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n476), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n466), .A2(new_n469), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n501), .A2(new_n513), .A3(new_n482), .ZN(new_n514));
  INV_X1    g313(.A(new_n497), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G183gat), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n470), .B1(new_n469), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n518), .A2(new_n449), .A3(new_n455), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n471), .A2(new_n473), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(new_n467), .A3(new_n470), .A4(new_n469), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n512), .A2(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G226gat), .A2(G233gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n445), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n522), .B2(KEYINPUT29), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n503), .A2(G226gat), .A3(G233gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n444), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT37), .ZN(new_n530));
  XOR2_X1   g329(.A(G8gat), .B(G36gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT78), .ZN(new_n532));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n529), .B2(KEYINPUT37), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT38), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n525), .A2(new_n528), .A3(new_n534), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n539), .A2(new_n537), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n431), .A2(new_n434), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n444), .B1(new_n390), .B2(new_n504), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(G228gat), .B2(G233gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n439), .A2(KEYINPUT83), .A3(new_n441), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n504), .B(new_n546), .C1(new_n444), .C2(KEYINPUT83), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n547), .A2(new_n389), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n374), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n444), .A2(new_n504), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n374), .B1(new_n550), .B2(new_n389), .ZN(new_n551));
  OAI211_X1 g350(.A(G228gat), .B(G233gat), .C1(new_n551), .C2(new_n544), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G50gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G78gat), .B(G106gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G22gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(new_n549), .B2(new_n552), .ZN(new_n560));
  OR3_X1    g359(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n556), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n423), .A2(KEYINPUT87), .A3(new_n424), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n379), .A2(new_n381), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n405), .A2(new_n400), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n383), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT39), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n426), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT39), .B1(new_n402), .B2(new_n403), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n571), .B(new_n573), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n417), .A2(KEYINPUT4), .ZN(new_n576));
  INV_X1    g375(.A(new_n381), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n568), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n570), .A3(new_n403), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n579), .B(new_n414), .C1(new_n569), .C2(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n572), .ZN(new_n581));
  INV_X1    g380(.A(new_n534), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n529), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT30), .A3(new_n539), .ZN(new_n584));
  OR3_X1    g383(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n582), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n575), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n563), .B1(new_n566), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n543), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n421), .A2(new_n426), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n433), .B1(new_n590), .B2(new_n415), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n563), .B1(new_n591), .B2(new_n586), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT84), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n512), .A2(new_n516), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n400), .A2(new_n594), .A3(new_n475), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n503), .A2(new_n395), .ZN(new_n596));
  AND2_X1   g395(.A1(G227gat), .A2(G233gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT74), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT32), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G15gat), .B(G43gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT75), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n216), .ZN(new_n608));
  INV_X1    g407(.A(G99gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT32), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(new_n600), .B2(new_n601), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT33), .B1(new_n600), .B2(new_n601), .ZN(new_n614));
  INV_X1    g413(.A(new_n610), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n597), .B1(new_n595), .B2(new_n596), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT77), .B(KEYINPUT34), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT34), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n611), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT36), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n611), .A2(new_n616), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n625), .B2(KEYINPUT76), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n627), .A3(new_n616), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n622), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n631));
  AOI221_X4 g430(.A(new_n612), .B1(new_n610), .B2(KEYINPUT33), .C1(new_n600), .C2(new_n601), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT36), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n592), .B(new_n593), .C1(new_n629), .C2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT76), .B1(new_n631), .B2(new_n632), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n628), .A3(new_n630), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n623), .A2(KEYINPUT36), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n623), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n561), .A2(new_n562), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n415), .A2(new_n590), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n434), .ZN(new_n644));
  INV_X1    g443(.A(new_n586), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT84), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n589), .A2(new_n635), .A3(new_n647), .ZN(new_n648));
  NOR4_X1   g447(.A1(new_n639), .A2(KEYINPUT35), .A3(new_n586), .A4(new_n563), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n432), .B1(new_n421), .B2(new_n426), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n564), .B2(new_n565), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(new_n651), .B2(new_n433), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n623), .A2(new_n561), .A3(new_n562), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n653), .A2(new_n637), .A3(new_n644), .A4(new_n645), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT35), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n214), .A2(new_n269), .A3(new_n270), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n212), .A2(new_n267), .A3(new_n213), .ZN(new_n659));
  NAND2_X1  g458(.A1(G229gat), .A2(G233gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT18), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT18), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n658), .A2(new_n663), .A3(new_n659), .A4(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n660), .B(KEYINPUT13), .Z(new_n666));
  INV_X1    g465(.A(new_n659), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n267), .B1(new_n212), .B2(new_n213), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT93), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT93), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G169gat), .B(G197gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT89), .B(KEYINPUT12), .Z(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n673), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n657), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT94), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT94), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n657), .A2(new_n688), .A3(new_n685), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n334), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n644), .A2(KEYINPUT106), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n644), .A2(KEYINPUT106), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT107), .B(G1gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1324gat));
  AOI21_X1  g495(.A(new_n211), .B1(new_n690), .B2(new_n586), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n688), .B1(new_n657), .B2(new_n685), .ZN(new_n698));
  INV_X1    g497(.A(new_n685), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT94), .B(new_n699), .C1(new_n648), .C2(new_n656), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT108), .B(KEYINPUT16), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G8gat), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n701), .A2(new_n645), .A3(new_n334), .A4(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n697), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT42), .B2(new_n704), .ZN(G1325gat));
  INV_X1    g505(.A(new_n639), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(G15gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n712));
  INV_X1    g511(.A(new_n641), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n709), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n711), .A2(new_n712), .B1(new_n690), .B2(new_n714), .ZN(G1326gat));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n687), .A2(new_n689), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  INV_X1    g518(.A(new_n334), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n563), .A4(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n563), .B(new_n720), .C1(new_n698), .C2(new_n700), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT110), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n721), .B2(new_n723), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n717), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n721), .A2(new_n723), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT111), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n716), .A3(new_n725), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1327gat));
  NOR2_X1   g531(.A1(new_n253), .A2(new_n332), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n305), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n698), .B2(new_n700), .ZN(new_n736));
  INV_X1    g535(.A(new_n693), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n736), .A2(G29gat), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT45), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n641), .A2(new_n646), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n651), .A2(new_n541), .A3(new_n433), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n566), .A2(new_n587), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n642), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n656), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n745), .B2(new_n304), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n304), .A2(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n648), .B2(new_n656), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n685), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n737), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n739), .A2(new_n753), .ZN(G1328gat));
  OR3_X1    g553(.A1(new_n736), .A2(G36gat), .A3(new_n645), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g555(.A(G36gat), .B1(new_n752), .B2(new_n645), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(KEYINPUT46), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(G1329gat));
  INV_X1    g558(.A(G43gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n736), .B2(new_n639), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n641), .A2(G43gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n752), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1330gat));
  NAND3_X1  g564(.A1(new_n718), .A2(KEYINPUT113), .A3(new_n735), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n736), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n642), .A2(G50gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  OAI21_X1  g570(.A(G50gat), .B1(new_n752), .B2(new_n642), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1331gat));
  AND4_X1   g575(.A1(new_n699), .A2(new_n307), .A3(new_n309), .A4(new_n332), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n745), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n737), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(new_n222), .ZN(G1332gat));
  AOI21_X1  g579(.A(new_n645), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT114), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n745), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n783), .B(new_n784), .Z(G1333gat));
  OAI21_X1  g584(.A(G71gat), .B1(new_n778), .B2(new_n713), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n707), .A2(new_n216), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g588(.A1(new_n778), .A2(new_n642), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n217), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n253), .A2(new_n685), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n592), .B1(new_n629), .B2(new_n634), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n543), .B2(new_n588), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n431), .A2(new_n434), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n795), .A2(new_n649), .B1(new_n654), .B2(KEYINPUT35), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n304), .B(new_n792), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n304), .A4(new_n792), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n333), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n272), .A3(new_n693), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n253), .A2(new_n685), .A3(new_n333), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n746), .A2(new_n748), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT115), .B1(new_n806), .B2(new_n737), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G85gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n806), .A2(KEYINPUT115), .A3(new_n737), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n802), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  AOI21_X1  g609(.A(new_n271), .B1(new_n805), .B2(new_n586), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n799), .A2(new_n800), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n333), .A2(G92gat), .A3(new_n645), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT52), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n812), .B2(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(new_n747), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n657), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n589), .A2(new_n740), .B1(new_n652), .B2(new_n655), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n305), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n819), .A2(new_n822), .A3(new_n586), .A4(new_n803), .ZN(new_n823));
  INV_X1    g622(.A(new_n271), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n817), .A2(KEYINPUT117), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n817), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n815), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n815), .C1(new_n826), .C2(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1337gat));
  OAI21_X1  g631(.A(G99gat), .B1(new_n806), .B2(new_n713), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n801), .A2(new_n609), .A3(new_n707), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1338gat));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  OAI21_X1  g635(.A(G106gat), .B1(new_n806), .B2(new_n642), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(G106gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n801), .A2(new_n840), .A3(new_n563), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n839), .B(new_n842), .ZN(G1339gat));
  NAND4_X1  g642(.A1(new_n307), .A2(new_n309), .A3(new_n699), .A4(new_n333), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n324), .A2(new_n846), .A3(new_n326), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n321), .B2(new_n322), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n318), .A2(G230gat), .A3(G233gat), .A4(new_n320), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n312), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT121), .B(KEYINPUT55), .C1(new_n847), .C2(new_n850), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n331), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n850), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT120), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n847), .A2(new_n850), .A3(new_n859), .A4(KEYINPUT55), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n660), .B1(new_n658), .B2(new_n659), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n667), .A2(new_n668), .A3(new_n666), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n679), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n684), .A2(new_n864), .ZN(new_n865));
  AND4_X1   g664(.A1(new_n304), .A2(new_n855), .A3(new_n861), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n332), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n858), .A2(new_n860), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n685), .A3(new_n331), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n853), .A2(new_n854), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n866), .B1(new_n305), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n844), .B1(new_n872), .B2(new_n253), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n639), .A2(new_n586), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n873), .A2(new_n642), .A3(new_n874), .A4(new_n693), .ZN(new_n875));
  INV_X1    g674(.A(G113gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(new_n699), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n873), .A2(new_n693), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n653), .A2(new_n637), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(new_n645), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n685), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(new_n876), .ZN(G1340gat));
  INV_X1    g683(.A(G120gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n875), .A2(new_n885), .A3(new_n333), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n882), .A2(new_n332), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n885), .ZN(G1341gat));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n338), .A3(new_n253), .ZN(new_n889));
  OAI21_X1  g688(.A(G127gat), .B1(new_n875), .B2(new_n308), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1342gat));
  NOR2_X1   g690(.A1(new_n305), .A2(new_n586), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n336), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n894));
  OAI21_X1  g693(.A(G134gat), .B1(new_n875), .B2(new_n305), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n641), .A2(new_n642), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n873), .A2(new_n645), .A3(new_n693), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n685), .A2(new_n355), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT55), .B1(new_n851), .B2(KEYINPUT122), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(KEYINPUT122), .B2(new_n851), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n861), .A3(new_n685), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n304), .B1(new_n906), .B2(new_n867), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n308), .B1(new_n907), .B2(new_n866), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n844), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n563), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n873), .A2(new_n912), .A3(new_n563), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n737), .A2(new_n586), .A3(new_n641), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n911), .A2(new_n685), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n903), .B1(new_n915), .B2(G141gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(G1344gat));
  INV_X1    g717(.A(new_n901), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n356), .A3(new_n332), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT57), .B(new_n642), .C1(new_n909), .C2(KEYINPUT124), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(KEYINPUT124), .B2(new_n909), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n873), .A2(new_n563), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n923), .A2(new_n332), .A3(new_n914), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT59), .B(new_n356), .C1(new_n928), .C2(new_n332), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n920), .B1(new_n927), .B2(new_n929), .ZN(G1345gat));
  NAND3_X1  g729(.A1(new_n919), .A2(new_n362), .A3(new_n253), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n928), .A2(new_n253), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n362), .ZN(G1346gat));
  NAND4_X1  g732(.A1(new_n878), .A2(new_n363), .A3(new_n892), .A4(new_n900), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n928), .A2(new_n304), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n363), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n693), .A2(new_n645), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n873), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(new_n880), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n685), .A3(new_n489), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n693), .A2(new_n645), .A3(new_n639), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n871), .A2(new_n305), .ZN(new_n942));
  INV_X1    g741(.A(new_n866), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n253), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n844), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n642), .B(new_n941), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n873), .A2(KEYINPUT125), .A3(new_n642), .A4(new_n941), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(new_n685), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n940), .B1(new_n451), .B2(new_n950), .ZN(G1348gat));
  NAND3_X1  g750(.A1(new_n939), .A2(new_n452), .A3(new_n332), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n948), .A2(new_n332), .A3(new_n949), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n452), .B2(new_n953), .ZN(G1349gat));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n517), .A3(new_n253), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n948), .A2(new_n253), .A3(new_n949), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n466), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n939), .A2(new_n469), .A3(new_n304), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n304), .A3(new_n949), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(G190gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n960), .B2(G190gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT61), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n960), .A2(G190gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n968), .B2(new_n962), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n959), .B1(new_n965), .B2(new_n969), .ZN(G1351gat));
  AND2_X1   g769(.A1(new_n938), .A2(new_n900), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n685), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n923), .A2(new_n925), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n693), .A2(new_n645), .A3(new_n641), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n685), .A2(G197gat), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1352gat));
  NAND3_X1  g776(.A1(new_n973), .A2(new_n332), .A3(new_n974), .ZN(new_n978));
  XOR2_X1   g777(.A(KEYINPUT127), .B(G204gat), .Z(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n333), .A2(new_n979), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n971), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g781(.A(new_n982), .B(KEYINPUT62), .Z(new_n983));
  NAND2_X1  g782(.A1(new_n980), .A2(new_n983), .ZN(G1353gat));
  NAND3_X1  g783(.A1(new_n971), .A2(new_n437), .A3(new_n253), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n923), .A2(new_n253), .A3(new_n925), .A4(new_n974), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n304), .A3(new_n974), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G218gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n971), .A2(new_n254), .A3(new_n304), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1355gat));
endmodule


