//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G50), .B2(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n209), .B(new_n225), .C1(new_n233), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT13), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G97), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G226), .A2(G1698), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n217), .B2(G1698), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n230), .A2(new_n262), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT69), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(G274), .C1(G41), .C2(G45), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT67), .B1(new_n269), .B2(new_n226), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n262), .A2(new_n271), .A3(G1), .A4(G13), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n270), .B2(new_n272), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n277), .B2(G238), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n254), .B1(new_n266), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n264), .A2(new_n254), .A3(new_n278), .A4(new_n265), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G169), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT14), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(KEYINPUT70), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n279), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G179), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(KEYINPUT14), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(G169), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n285), .A2(new_n287), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n228), .A2(new_n229), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n255), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n297), .A2(new_n298), .B1(new_n232), .B2(G68), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n202), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n221), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT12), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n295), .B1(new_n267), .B2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G68), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT71), .Z(new_n312));
  OR2_X1    g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n203), .A2(G20), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n315), .B1(new_n316), .B2(new_n301), .C1(new_n297), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n295), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n306), .A2(new_n202), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n310), .A2(G50), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G222), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n260), .A2(G1698), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT68), .ZN(new_n331));
  INV_X1    g0131(.A(G223), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n329), .B1(new_n298), .B2(new_n260), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n263), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n273), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n277), .A2(G226), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n323), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G179), .B2(new_n338), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(new_n322), .B(KEYINPUT9), .Z(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n338), .B2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n344), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n342), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n328), .A2(G232), .B1(G107), .B2(new_n327), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n331), .B2(new_n222), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n334), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n277), .A2(G244), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n354), .A2(new_n336), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT15), .B(G87), .Z(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n297), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n317), .A2(new_n301), .B1(new_n232), .B2(new_n298), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n295), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n306), .A2(new_n298), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n310), .A2(G77), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n354), .A2(new_n336), .A3(new_n355), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n339), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n358), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n314), .A2(new_n351), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n313), .B1(new_n289), .B2(G190), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n282), .A2(G200), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n255), .A2(KEYINPUT73), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G33), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT3), .ZN(new_n379));
  INV_X1    g0179(.A(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n332), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(G226), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n379), .A2(new_n325), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n273), .B1(new_n385), .B2(new_n334), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n217), .B(new_n276), .C1(new_n270), .C2(new_n272), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(G200), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n263), .B1(new_n383), .B2(new_n384), .ZN(new_n390));
  NOR4_X1   g0190(.A1(new_n390), .A2(new_n387), .A3(G190), .A4(new_n273), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n375), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n385), .A2(new_n334), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n393), .A2(new_n345), .A3(new_n336), .A4(new_n388), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n390), .A2(new_n273), .A3(new_n387), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(KEYINPUT74), .C1(new_n395), .C2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(G58), .B(G68), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(G20), .B1(G159), .B2(new_n300), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n379), .B2(new_n325), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n325), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT73), .B(G33), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n405), .A2(KEYINPUT7), .A3(G20), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT16), .B(new_n399), .C1(new_n402), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n401), .A2(G20), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT3), .B1(new_n376), .B2(new_n378), .ZN(new_n410));
  INV_X1    g0210(.A(new_n326), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n401), .B1(new_n260), .B2(G20), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n221), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n399), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n416), .A3(new_n295), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n317), .A2(new_n305), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n310), .B2(new_n317), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n397), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n417), .A2(new_n419), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n392), .B2(new_n396), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n395), .A2(G179), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n339), .B2(new_n395), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n354), .A2(G190), .A3(new_n336), .A4(new_n355), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n367), .B(new_n435), .C1(new_n356), .C2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n374), .A2(new_n427), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n371), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n379), .A2(G244), .A3(new_n380), .A4(new_n325), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT4), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n325), .A2(new_n326), .A3(G250), .A4(G1698), .ZN(new_n443));
  AND2_X1   g0243(.A1(KEYINPUT4), .A2(G244), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n325), .A2(new_n326), .A3(new_n444), .A4(new_n380), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n263), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT5), .B(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n275), .A2(G1), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n270), .A2(new_n272), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G257), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n449), .A2(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n273), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G169), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n451), .A2(G257), .B1(new_n273), .B2(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n441), .B2(new_n440), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(G179), .C1(new_n459), .C2(new_n263), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n218), .B1(new_n412), .B2(new_n413), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n462), .A2(new_n256), .A3(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n465), .A2(new_n232), .B1(new_n298), .B2(new_n301), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n295), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n305), .A2(G97), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n255), .A2(G1), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n295), .A2(new_n306), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G97), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n456), .A2(new_n460), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n213), .A2(new_n380), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n380), .A2(G257), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n379), .A2(new_n325), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G294), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(new_n404), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n334), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n451), .A2(G264), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n454), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n478), .A2(new_n334), .B1(G264), .B2(new_n451), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G190), .A3(new_n454), .ZN(new_n484));
  INV_X1    g0284(.A(new_n295), .ZN(new_n485));
  INV_X1    g0285(.A(new_n469), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(G107), .A3(new_n305), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(KEYINPUT25), .C1(new_n305), .C2(G107), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n489), .A2(KEYINPUT25), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(KEYINPUT25), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n306), .A2(new_n491), .A3(new_n218), .A4(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n487), .A2(new_n488), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  NOR4_X1   g0294(.A1(new_n295), .A2(new_n306), .A3(new_n218), .A4(new_n469), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n490), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT83), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n376), .B2(new_n378), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n232), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n232), .A2(G87), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n327), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n218), .A2(G20), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n504), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n379), .A2(KEYINPUT22), .A3(new_n325), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n499), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n260), .A2(new_n510), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n503), .B1(new_n501), .B2(new_n232), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT24), .A3(new_n511), .A4(new_n508), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n295), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n482), .A2(new_n484), .A3(new_n498), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT75), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n467), .A2(new_n471), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n467), .B2(new_n471), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n457), .B1(new_n459), .B2(new_n263), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n521), .A2(new_n522), .B1(new_n345), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(G200), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT76), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT76), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n527), .B(G200), .C1(new_n448), .C2(new_n455), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n473), .B(new_n518), .C1(new_n524), .C2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n405), .A2(KEYINPUT78), .A3(G244), .A4(G1698), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n379), .A2(G244), .A3(G1698), .A4(new_n325), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT78), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n501), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n405), .A2(KEYINPUT77), .A3(G238), .A4(new_n380), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n379), .A2(G238), .A3(new_n380), .A4(new_n325), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT77), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n334), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n270), .A2(new_n272), .ZN(new_n543));
  OR3_X1    g0343(.A1(new_n275), .A2(G1), .A3(G274), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(G250), .C2(new_n450), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n405), .A2(new_n232), .A3(G68), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n297), .B2(new_n256), .ZN(new_n550));
  NOR3_X1   g0350(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(new_n257), .B2(KEYINPUT19), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n548), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n295), .B1(new_n306), .B2(new_n360), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n470), .A2(G87), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n542), .A2(G190), .A3(new_n545), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n547), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n546), .A2(new_n339), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n542), .A2(new_n357), .A3(new_n545), .ZN(new_n560));
  INV_X1    g0360(.A(new_n470), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n554), .B1(new_n360), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n530), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  INV_X1    g0366(.A(G303), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n325), .B2(new_n326), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G257), .A2(G1698), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n219), .B2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n405), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n571), .B2(new_n263), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n451), .A2(G270), .B1(new_n273), .B2(new_n453), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n379), .A3(new_n325), .ZN(new_n574));
  INV_X1    g0374(.A(new_n568), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n334), .A3(KEYINPUT79), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT80), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT80), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n572), .A2(new_n580), .A3(new_n573), .A4(new_n577), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(G190), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n500), .A2(G20), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n446), .B(new_n232), .C1(G33), .C2(new_n256), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n295), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n295), .A2(KEYINPUT20), .A3(new_n585), .A4(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n470), .A2(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n306), .A2(new_n500), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n583), .A2(new_n584), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT81), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n583), .A2(new_n598), .A3(new_n584), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(G169), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT21), .B1(new_n582), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n604), .B(new_n601), .C1(new_n579), .C2(new_n581), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n572), .A2(G179), .A3(new_n573), .A4(new_n577), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n595), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n517), .A2(new_n498), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n481), .A2(new_n339), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n483), .A2(new_n357), .A3(new_n454), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NOR4_X1   g0411(.A1(new_n603), .A2(new_n605), .A3(new_n607), .A4(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n439), .A2(new_n565), .A3(new_n600), .A4(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n313), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n283), .B(new_n291), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n290), .A2(new_n287), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n370), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n427), .B(new_n374), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n434), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n348), .A2(new_n350), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n342), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n409), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n377), .A2(G33), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n255), .A2(KEYINPUT73), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n324), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n626), .B2(new_n326), .ZN(new_n627));
  INV_X1    g0427(.A(new_n413), .ZN(new_n628));
  OAI21_X1  g0428(.A(G107), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n464), .A2(new_n462), .ZN(new_n630));
  INV_X1    g0430(.A(new_n463), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(G20), .B1(G77), .B2(new_n300), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n485), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n471), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT75), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n456), .A2(new_n460), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n520), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT84), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT84), .A4(new_n520), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n558), .A3(new_n563), .A4(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n564), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .A3(new_n472), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n642), .A2(KEYINPUT85), .A3(new_n643), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n563), .ZN(new_n651));
  INV_X1    g0451(.A(new_n603), .ZN(new_n652));
  INV_X1    g0452(.A(new_n607), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n582), .A2(KEYINPUT21), .A3(new_n602), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n565), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n439), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n622), .A2(new_n659), .ZN(G369));
  NOR2_X1   g0460(.A1(new_n603), .A2(new_n605), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n653), .ZN(new_n662));
  INV_X1    g0462(.A(G13), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n267), .ZN(new_n665));
  XNOR2_X1  g0465(.A(KEYINPUT86), .B(KEYINPUT27), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n594), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n600), .A2(new_n672), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n662), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n676));
  XOR2_X1   g0476(.A(KEYINPUT88), .B(G330), .Z(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(KEYINPUT87), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n655), .A2(new_n671), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n608), .A2(new_n671), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n518), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n655), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n676), .A2(new_n677), .A3(new_n678), .A4(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n679), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n671), .B1(new_n661), .B2(new_n653), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n207), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G1), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n551), .A2(new_n500), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n234), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(new_n671), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n600), .A2(new_n612), .A3(new_n565), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n542), .A2(new_n483), .A3(new_n545), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT90), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n542), .A2(new_n483), .A3(new_n699), .A4(new_n545), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n606), .A2(new_n523), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n582), .A2(new_n523), .A3(new_n546), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n481), .A2(new_n357), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n706), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n701), .A2(new_n711), .A3(new_n704), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n671), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n696), .A2(new_n714), .A3(KEYINPUT31), .ZN(new_n715));
  XNOR2_X1  g0515(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(new_n671), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n677), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n671), .B1(new_n650), .B2(new_n657), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n523), .A2(new_n345), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n636), .B2(new_n520), .ZN(new_n724));
  INV_X1    g0524(.A(new_n528), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n527), .B1(new_n523), .B2(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n472), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n518), .A3(new_n563), .A4(new_n558), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT93), .B1(new_n612), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT93), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n565), .A2(new_n731), .A3(new_n656), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n563), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n642), .A2(new_n734), .A3(new_n643), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n642), .A2(new_n643), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n558), .A2(new_n563), .A3(new_n472), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n643), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT29), .B(new_n695), .C1(new_n733), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n720), .B1(new_n722), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n694), .B1(new_n742), .B2(G1), .ZN(G364));
  NAND2_X1  g0543(.A1(new_n676), .A2(new_n678), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n677), .ZN(new_n746));
  INV_X1    g0546(.A(new_n677), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n691), .B1(G45), .B2(new_n664), .ZN(new_n749));
  OR3_X1    g0549(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n232), .A2(new_n357), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G190), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n436), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G326), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n751), .A2(new_n345), .A3(G200), .ZN(new_n760));
  OR2_X1    g0560(.A1(KEYINPUT33), .A2(G317), .ZN(new_n761));
  NAND2_X1  g0561(.A1(KEYINPUT33), .A2(G317), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n436), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n232), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n751), .A2(new_n345), .A3(new_n436), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n327), .B1(new_n766), .B2(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n232), .B1(new_n771), .B2(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n763), .B(new_n770), .C1(G294), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n764), .A2(G20), .A3(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G303), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n752), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n765), .A2(new_n771), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(G322), .B1(G329), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n759), .A2(new_n774), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n260), .B1(new_n775), .B2(new_n212), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n256), .ZN(new_n789));
  INV_X1    g0589(.A(new_n768), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n785), .B(new_n789), .C1(G77), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n766), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n758), .A2(G50), .B1(G107), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  OAI21_X1  g0594(.A(KEYINPUT32), .B1(new_n779), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n778), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n221), .B2(new_n760), .C1(new_n796), .C2(new_n216), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(KEYINPUT96), .B2(new_n784), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n791), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n779), .A2(KEYINPUT32), .A3(new_n794), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n782), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n231), .B1(G20), .B2(new_n339), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT94), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n260), .A2(G355), .A3(new_n207), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n249), .A2(new_n275), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n405), .A2(new_n688), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G45), .B2(new_n235), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(G116), .B2(new_n207), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n801), .A2(new_n802), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n805), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n749), .B(new_n813), .C1(new_n745), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n750), .A2(new_n815), .ZN(G396));
  INV_X1    g0616(.A(new_n721), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n366), .A2(new_n671), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n437), .A2(new_n818), .B1(new_n369), .B2(new_n358), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n358), .A2(new_n369), .A3(new_n695), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT99), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT99), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n366), .B1(new_n368), .B2(G200), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(new_n435), .B1(new_n366), .B2(new_n671), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n820), .C1(new_n618), .C2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n817), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT100), .B1(new_n721), .B2(new_n827), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n832), .A2(new_n719), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n720), .B1(new_n835), .B2(new_n831), .ZN(new_n836));
  INV_X1    g0636(.A(new_n749), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n802), .A2(new_n803), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n298), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n827), .B2(new_n804), .ZN(new_n841));
  INV_X1    g0641(.A(new_n760), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G143), .A2(new_n778), .B1(new_n842), .B2(G150), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n794), .B2(new_n768), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n758), .B2(G137), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT34), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n773), .A2(G58), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n776), .A2(G50), .B1(new_n792), .B2(G68), .ZN(new_n848));
  INV_X1    g0648(.A(new_n405), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G132), .B2(new_n780), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n757), .A2(new_n567), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n792), .A2(G87), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n769), .B2(new_n779), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n789), .B(new_n852), .C1(KEYINPUT98), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n776), .A2(G107), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(KEYINPUT98), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n260), .B(new_n857), .C1(G294), .C2(new_n778), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G116), .A2(new_n790), .B1(new_n842), .B2(G283), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n855), .A2(new_n856), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n837), .B(new_n841), .C1(new_n802), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n838), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  INV_X1    g0664(.A(KEYINPUT108), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n701), .A2(new_n704), .A3(new_n711), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n711), .B1(new_n701), .B2(new_n704), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n708), .A2(new_n709), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n869), .B2(new_n695), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n713), .A2(KEYINPUT108), .A3(new_n671), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n717), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n696), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n828), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n293), .A2(new_n313), .A3(new_n695), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n372), .A2(new_n373), .B1(new_n313), .B2(new_n671), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n617), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n669), .B(KEYINPUT102), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n424), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(KEYINPUT103), .B(new_n885), .C1(new_n417), .C2(new_n419), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n421), .B(new_n430), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n890));
  INV_X1    g0690(.A(new_n887), .ZN(new_n891));
  INV_X1    g0691(.A(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n424), .A2(new_n429), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n425), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT104), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n893), .B2(new_n895), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n893), .B1(new_n427), .B2(new_n434), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n882), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n399), .B1(new_n402), .B2(new_n406), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n408), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n407), .A2(new_n295), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n419), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n669), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n908), .B1(new_n429), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n421), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n890), .A2(new_n897), .B1(KEYINPUT37), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n434), .A2(new_n423), .A3(new_n426), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n909), .A3(new_n908), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT40), .B1(new_n904), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n880), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n920));
  NAND2_X1  g0720(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n898), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n917), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n880), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n872), .A2(new_n874), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n439), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n926), .B(new_n928), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n677), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n741), .B(new_n439), .C1(KEYINPUT29), .C2(new_n721), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n622), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n922), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n899), .B1(new_n890), .B2(new_n897), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n881), .B1(new_n936), .B2(new_n902), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT39), .B1(new_n923), .B2(new_n917), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n934), .A2(new_n937), .A3(new_n941), .A4(new_n935), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n876), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n434), .A2(new_n886), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n820), .B(KEYINPUT101), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n721), .B2(new_n827), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n878), .ZN(new_n949));
  INV_X1    g0749(.A(new_n924), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n933), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n267), .B2(new_n664), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n500), .B1(new_n632), .B2(KEYINPUT35), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(new_n233), .C1(KEYINPUT35), .C2(new_n632), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  OAI21_X1  g0757(.A(G77), .B1(new_n216), .B2(new_n221), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n958), .A2(new_n234), .B1(G50), .B2(new_n221), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(G1), .A3(new_n663), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(new_n957), .A3(new_n960), .ZN(G367));
  NAND2_X1  g0761(.A1(new_n686), .A2(new_n684), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n636), .A2(new_n520), .A3(new_n671), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n728), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n638), .B2(new_n695), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n962), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(new_n966), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n683), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n685), .B(new_n682), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n748), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n742), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT110), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n689), .B(KEYINPUT41), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n742), .ZN(new_n981));
  INV_X1    g0781(.A(new_n975), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n748), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n981), .B1(new_n983), .B2(new_n973), .ZN(new_n984));
  INV_X1    g0784(.A(new_n979), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT110), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n267), .B1(new_n664), .B2(G45), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n980), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n685), .A2(new_n728), .A3(new_n682), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT42), .Z(new_n990));
  AOI21_X1  g0790(.A(new_n472), .B1(new_n965), .B2(new_n611), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n671), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n556), .A2(new_n695), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n647), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n563), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n683), .A2(new_n966), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n988), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(G143), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n757), .A2(new_n1004), .B1(new_n202), .B2(new_n768), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G159), .B2(new_n842), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n788), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(G68), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT112), .B(G137), .Z(new_n1009));
  OAI22_X1  g0809(.A1(new_n779), .A2(new_n1009), .B1(new_n775), .B2(new_n216), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G150), .B2(new_n778), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n792), .A2(G77), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n260), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT111), .Z(new_n1014));
  NAND4_X1  g0814(.A1(new_n1006), .A2(new_n1008), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n757), .A2(new_n769), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n766), .A2(new_n256), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n776), .A2(G116), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT46), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n796), .A2(new_n567), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(new_n1019), .C2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(G317), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1022), .A2(new_n779), .B1(new_n772), .B2(new_n218), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n405), .B(new_n1023), .C1(G283), .C2(new_n790), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(new_n477), .C2(new_n760), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1015), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n802), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n994), .A2(new_n805), .A3(new_n995), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n810), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n807), .B1(new_n207), .B2(new_n360), .C1(new_n244), .C2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n749), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1003), .A2(new_n1032), .ZN(G387));
  OR3_X1    g0833(.A1(new_n983), .A2(KEYINPUT115), .A3(new_n742), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT115), .B1(new_n983), .B2(new_n742), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n983), .A2(new_n742), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n689), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n987), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n983), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n405), .B1(new_n317), .B2(new_n760), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1007), .A2(new_n359), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n202), .B2(new_n796), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT113), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(G77), .C2(new_n776), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n758), .A2(G159), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n780), .A2(G150), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1017), .B1(G68), .B2(new_n790), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n775), .A2(new_n477), .B1(new_n772), .B2(new_n767), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G317), .A2(new_n778), .B1(new_n842), .B2(G311), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n567), .B2(new_n768), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n758), .B2(G322), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1052), .B2(KEYINPUT48), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT114), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(KEYINPUT48), .B2(new_n1052), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT49), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n780), .A2(G326), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n849), .B(new_n1057), .C1(new_n500), .C2(new_n766), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1048), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n802), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n682), .A2(new_n814), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n810), .B1(new_n241), .B2(new_n275), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n692), .A2(new_n207), .A3(new_n260), .ZN(new_n1063));
  AOI211_X1 g0863(.A(G45), .B(new_n692), .C1(G68), .C2(G77), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n317), .A2(G50), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT50), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1062), .A2(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n207), .A2(G107), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n807), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1060), .A2(new_n749), .A3(new_n1061), .A4(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1037), .A2(new_n1039), .A3(new_n1070), .ZN(G393));
  AOI21_X1  g0871(.A(new_n690), .B1(new_n1036), .B2(new_n974), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n974), .B2(new_n1036), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n966), .A2(new_n805), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n758), .A2(G150), .B1(G159), .B2(new_n778), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1075), .A2(KEYINPUT51), .B1(new_n1004), .B2(new_n779), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(KEYINPUT51), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n849), .B1(G50), .B2(new_n842), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n317), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(new_n790), .B1(new_n776), .B2(G68), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n853), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1076), .B(new_n1081), .C1(G77), .C2(new_n1007), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n757), .A2(new_n1022), .B1(new_n769), .B2(new_n796), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n790), .A2(G294), .B1(new_n773), .B2(G116), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n775), .A2(new_n767), .B1(new_n766), .B2(new_n218), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n260), .B(new_n1086), .C1(G322), .C2(new_n780), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G303), .B2(new_n842), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n802), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n807), .B1(new_n256), .B2(new_n207), .C1(new_n252), .C2(new_n1030), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1074), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n973), .A2(new_n1038), .B1(new_n749), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1073), .A2(new_n1093), .ZN(G390));
  OAI211_X1 g0894(.A(new_n695), .B(new_n827), .C1(new_n733), .C2(new_n740), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n820), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n617), .A2(new_n877), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n944), .B1(new_n934), .B2(new_n937), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1097), .B1(new_n1095), .B2(new_n820), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n876), .B1(new_n904), .B2(new_n917), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT116), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n876), .B1(new_n948), .B2(new_n878), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1107), .A2(new_n940), .A3(new_n939), .A4(new_n942), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n715), .A2(new_n677), .A3(new_n718), .A4(new_n827), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n879), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1106), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n875), .A2(G330), .A3(new_n879), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n820), .B(new_n1095), .C1(new_n1109), .C2(new_n878), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n927), .A2(G330), .A3(new_n827), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n878), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n879), .B1(new_n875), .B2(G330), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT117), .B1(new_n1121), .B2(new_n1115), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1113), .B1(new_n1110), .B2(new_n879), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n948), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1120), .A2(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n927), .A2(new_n439), .A3(G330), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n932), .A2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1112), .A2(new_n1114), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1100), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1103), .A2(new_n1104), .A3(KEYINPUT116), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1108), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1113), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1108), .B(new_n1111), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1128), .A2(new_n1138), .A3(new_n689), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n803), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n775), .A2(new_n316), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1143), .A2(KEYINPUT53), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(KEYINPUT53), .B1(new_n778), .B2(G132), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n792), .A2(G50), .B1(new_n780), .B2(G125), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n260), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n758), .A2(G128), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n760), .B2(new_n1009), .C1(new_n794), .C2(new_n788), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT54), .B(G143), .Z(new_n1150));
  AOI211_X1 g0950(.A(new_n1147), .B(new_n1149), .C1(new_n790), .C2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n792), .A2(G68), .B1(new_n780), .B2(G294), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1152), .B(new_n327), .C1(new_n212), .C2(new_n775), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1007), .A2(G77), .B1(G97), .B2(new_n790), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n218), .B2(new_n760), .C1(new_n757), .C2(new_n767), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(G116), .C2(new_n778), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n802), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n839), .A2(new_n317), .ZN(new_n1158));
  AND4_X1   g0958(.A1(new_n749), .A2(new_n1141), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1160), .B2(new_n1038), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1139), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT118), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1139), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(G378));
  AOI21_X1  g0966(.A(G41), .B1(new_n758), .B2(G116), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(new_n849), .C1(new_n218), .C2(new_n796), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n766), .A2(new_n216), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G77), .B2(new_n776), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1008), .A2(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n256), .B2(new_n760), .C1(new_n767), .C2(new_n779), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1168), .B(new_n1172), .C1(new_n359), .C2(new_n790), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT58), .Z(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n625), .B2(KEYINPUT3), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n758), .A2(G125), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G132), .A2(new_n842), .B1(new_n790), .B2(G137), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT119), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1150), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1178), .B1(new_n316), .B2(new_n788), .C1(new_n775), .C2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1176), .B(new_n1180), .C1(G128), .C2(new_n778), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT59), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G33), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G41), .B1(new_n780), .B2(G124), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n794), .C2(new_n766), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1174), .B1(G50), .B2(new_n1175), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT120), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n802), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n839), .A2(new_n202), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n323), .A2(new_n669), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n351), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n803), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1189), .A2(new_n749), .A3(new_n1190), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n919), .A2(G330), .A3(new_n925), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1194), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n945), .A2(new_n951), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n945), .B2(new_n951), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n952), .A2(new_n1194), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n945), .A2(new_n951), .A3(new_n1199), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1202), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1197), .B1(new_n1207), .B2(new_n1038), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1127), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1140), .A2(new_n1107), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1137), .B1(new_n1211), .B2(new_n1113), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1119), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1121), .A2(new_n1115), .A3(KEYINPUT117), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1130), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1210), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1207), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n690), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1207), .A2(new_n1217), .A3(KEYINPUT57), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1209), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1216), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n985), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT121), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n878), .A2(new_n803), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n796), .A2(new_n1009), .B1(new_n760), .B2(new_n1179), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n758), .B2(G132), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT122), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n776), .A2(G159), .B1(new_n780), .B2(G128), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1169), .B(new_n849), .C1(G150), .C2(new_n790), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G50), .B2(new_n1007), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n260), .B1(new_n758), .B2(G294), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n842), .A2(G116), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1012), .A3(new_n1041), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n779), .A2(new_n567), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n775), .A2(new_n256), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n796), .A2(new_n767), .B1(new_n218), .B2(new_n768), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n802), .B1(new_n1235), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n839), .A2(new_n221), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1228), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1215), .A2(new_n1038), .B1(new_n749), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1227), .A2(new_n1246), .ZN(G381));
  INV_X1    g1047(.A(G390), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1003), .A3(new_n1032), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1249), .A2(G396), .A3(G393), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1162), .A2(KEYINPUT123), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1139), .A2(new_n1161), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1222), .A2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G381), .A2(G384), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1250), .A2(new_n1255), .A3(new_n1256), .ZN(G407));
  INV_X1    g1057(.A(G213), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1255), .B2(new_n670), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(G407), .ZN(G409));
  INV_X1    g1060(.A(G396), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(G393), .B(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1248), .A2(new_n1003), .A3(new_n1032), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1248), .B1(new_n1003), .B2(new_n1032), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G387), .A2(G390), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(G396), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1249), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1258), .A2(G343), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G2897), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1225), .A2(KEYINPUT60), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1224), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n689), .A3(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1275), .A2(G384), .A3(new_n1246), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1275), .B2(new_n1246), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1246), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n863), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(G384), .A3(new_n1246), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1271), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1208), .B1(new_n985), .B2(new_n1218), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1222), .A2(G378), .B1(new_n1254), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1286), .B2(new_n1270), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1222), .A2(G378), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1254), .A2(new_n1285), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1270), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1287), .A2(new_n1288), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1270), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1288), .A3(new_n1296), .A4(new_n1293), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1269), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1296), .A4(new_n1293), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT127), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1276), .A2(new_n1277), .A3(new_n1271), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1282), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1278), .A2(new_n1283), .A3(KEYINPUT126), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1306), .B(new_n1307), .C1(new_n1270), .C2(new_n1286), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1269), .A2(KEYINPUT61), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1291), .A2(new_n1310), .A3(KEYINPUT63), .A4(new_n1293), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1302), .A2(new_n1308), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1286), .A2(new_n1270), .A3(new_n1292), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1295), .A2(new_n1296), .A3(new_n1293), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1315), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(KEYINPUT125), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1300), .B1(new_n1312), .B2(new_n1320), .ZN(G405));
  NAND2_X1  g1121(.A1(G375), .A2(new_n1254), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1269), .A2(new_n1289), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1289), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1292), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1323), .A2(new_n1293), .A3(new_n1325), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


