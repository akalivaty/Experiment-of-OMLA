//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  XOR2_X1   g000(.A(KEYINPUT24), .B(G110), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n193), .B1(new_n190), .B2(new_n192), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n188), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n191), .A2(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(new_n198), .B2(KEYINPUT77), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT77), .B1(new_n189), .B2(G119), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n202), .A3(new_n192), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n197), .B1(G110), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT78), .B1(new_n206), .B2(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT16), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(new_n212), .A3(new_n205), .A4(G125), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n207), .A2(new_n210), .A3(G146), .A4(new_n213), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n204), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n192), .B1(new_n200), .B2(new_n201), .ZN(new_n221));
  AOI211_X1 g035(.A(KEYINPUT77), .B(KEYINPUT23), .C1(new_n189), .C2(G119), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(G110), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n189), .A2(G119), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT76), .B1(new_n198), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n187), .B1(new_n225), .B2(new_n194), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT79), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n188), .B1(new_n195), .B2(new_n196), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n229));
  INV_X1    g043(.A(G110), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n199), .A2(new_n202), .A3(new_n230), .A4(new_n192), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n206), .A2(new_n209), .A3(new_n215), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT80), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT80), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n206), .A2(new_n209), .A3(new_n236), .A4(new_n215), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n217), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n220), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  AOI211_X1 g055(.A(KEYINPUT81), .B(new_n239), .C1(new_n227), .C2(new_n232), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n219), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT82), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n219), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT22), .B(G137), .ZN(new_n247));
  INV_X1    g061(.A(G953), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n247), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n244), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n233), .A2(new_n240), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT81), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n233), .A2(new_n220), .A3(new_n240), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n255), .A2(new_n256), .B1(new_n218), .B2(new_n204), .ZN(new_n257));
  AOI21_X1  g071(.A(G902), .B1(new_n257), .B2(new_n250), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n252), .B2(new_n258), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n262));
  INV_X1    g076(.A(G234), .ZN(new_n263));
  OAI21_X1  g077(.A(G217), .B1(new_n263), .B2(G902), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT75), .ZN(new_n265));
  NOR4_X1   g079(.A1(new_n260), .A2(new_n261), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n252), .A2(new_n258), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n267), .B2(KEYINPUT25), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT83), .B1(new_n268), .B2(new_n259), .ZN(new_n269));
  INV_X1    g083(.A(new_n252), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n243), .A2(new_n251), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n265), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n266), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT2), .B(G113), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n191), .A2(G116), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G119), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n279), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  INV_X1    g103(.A(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G137), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT11), .ZN(new_n292));
  INV_X1    g106(.A(G137), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(G134), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n290), .A2(KEYINPUT11), .A3(G137), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n289), .B(new_n291), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT65), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT11), .B1(new_n290), .B2(G137), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n293), .A3(G134), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n298), .A2(new_n299), .B1(new_n290), .B2(G137), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n289), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n215), .A2(G143), .ZN(new_n304));
  INV_X1    g118(.A(G143), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n305), .A2(KEYINPUT64), .A3(G146), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT64), .B1(new_n305), .B2(G146), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(G143), .B2(new_n215), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n311), .B(KEYINPUT1), .C1(new_n305), .C2(G146), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G128), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n305), .A2(G146), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n304), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G143), .B(G146), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT68), .A3(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n290), .B2(G137), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n303), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT0), .A2(G128), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT0), .A2(G128), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n308), .A2(new_n333), .B1(new_n321), .B2(new_n331), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n300), .B2(new_n289), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT66), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n340), .B2(new_n303), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n288), .B1(new_n329), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n303), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n334), .ZN(new_n344));
  INV_X1    g158(.A(new_n288), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n303), .A2(new_n324), .A3(new_n328), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n278), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n329), .A2(new_n341), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT28), .B1(new_n349), .B2(new_n345), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G101), .ZN(new_n352));
  INV_X1    g166(.A(G237), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n248), .A3(G210), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n352), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT30), .B1(new_n329), .B2(new_n341), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n344), .A2(new_n363), .A3(new_n346), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n345), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n347), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n358), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n347), .A2(new_n278), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n357), .B(KEYINPUT71), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n342), .A2(new_n347), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n278), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n359), .B(new_n367), .C1(new_n371), .C2(KEYINPUT74), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n371), .A2(KEYINPUT74), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n361), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G472), .ZN(new_n375));
  INV_X1    g189(.A(new_n369), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n348), .B2(new_n350), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT72), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(new_n376), .C1(new_n348), .C2(new_n350), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n362), .A2(new_n364), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n366), .B1(new_n381), .B2(new_n288), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT31), .B1(new_n382), .B2(new_n357), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT31), .ZN(new_n384));
  NOR4_X1   g198(.A1(new_n365), .A2(new_n384), .A3(new_n366), .A4(new_n358), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n378), .B(new_n380), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT32), .ZN(new_n387));
  NOR2_X1   g201(.A1(G472), .A2(G902), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n388), .B(KEYINPUT73), .Z(new_n389));
  AND3_X1   g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n375), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT9), .B(G234), .ZN(new_n393));
  OAI21_X1  g207(.A(G221), .B1(new_n393), .B2(G902), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT84), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT12), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G104), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(G107), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n397), .A2(G107), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n400), .A2(G104), .ZN(new_n406));
  OAI21_X1  g220(.A(G101), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n315), .A2(new_n323), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT68), .B1(new_n321), .B2(new_n316), .ZN(new_n412));
  AND4_X1   g226(.A1(KEYINPUT68), .A2(new_n316), .A3(new_n304), .A4(new_n317), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n310), .A2(new_n189), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(new_n321), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT85), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n409), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n343), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n396), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n416), .B1(new_n323), .B2(new_n411), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n408), .B1(new_n423), .B2(new_n418), .ZN(new_n424));
  OAI211_X1 g238(.A(KEYINPUT12), .B(new_n343), .C1(new_n424), .C2(new_n409), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n248), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G101), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT4), .A3(new_n404), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n433), .A3(G101), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n334), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n315), .A2(new_n323), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n419), .A2(new_n410), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n429), .B1(new_n441), .B2(new_n421), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n426), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT86), .B1(new_n422), .B2(new_n425), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT87), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n442), .A4(new_n426), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n441), .A2(new_n421), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n441), .A2(new_n421), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n429), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G469), .ZN(new_n454));
  INV_X1    g268(.A(G902), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n422), .A2(new_n425), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n450), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n459), .A2(new_n429), .B1(new_n449), .B2(new_n442), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(G469), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n395), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n436), .A2(new_n208), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n335), .A2(G125), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n465), .B2(new_n466), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n432), .A2(new_n288), .A3(new_n434), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n284), .A2(KEYINPUT5), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g291(.A(G113), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n476), .A2(new_n479), .B1(new_n284), .B2(new_n280), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n410), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n474), .B1(new_n482), .B2(KEYINPUT89), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n475), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n475), .A2(new_n481), .A3(new_n474), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT6), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n473), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n472), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n467), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n410), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n496), .A2(new_n480), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n474), .B(KEYINPUT8), .Z(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n496), .B2(new_n480), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n465), .A2(KEYINPUT7), .A3(new_n471), .A4(new_n466), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n487), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n455), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n464), .B1(new_n491), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n500), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT7), .B1(new_n465), .B2(new_n466), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n506), .A2(new_n472), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n503), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n490), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n483), .A2(new_n485), .B1(KEYINPUT6), .B2(new_n487), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n511), .A2(new_n512), .B1(new_n470), .B2(new_n472), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n513), .A3(new_n463), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n514), .A3(KEYINPUT91), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n463), .B1(new_n510), .B2(new_n513), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT88), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n353), .A2(new_n248), .A3(G214), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(KEYINPUT92), .B2(new_n305), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT92), .B(G143), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G131), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n523), .B(new_n289), .C1(new_n522), .C2(new_n524), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n524), .A2(new_n522), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n289), .B1(new_n530), .B2(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n529), .A2(new_n532), .A3(new_n217), .A4(new_n216), .ZN(new_n533));
  XNOR2_X1  g347(.A(G113), .B(G122), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(new_n397), .ZN(new_n535));
  AND2_X1   g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n525), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n536), .A3(new_n523), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n215), .B1(new_n206), .B2(new_n209), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT93), .B1(new_n238), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n544), .B(new_n541), .C1(new_n235), .C2(new_n237), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n540), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n533), .A2(new_n535), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n535), .B1(new_n533), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(KEYINPUT95), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n455), .ZN(new_n553));
  OAI21_X1  g367(.A(G475), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(G475), .A2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n557));
  XNOR2_X1  g371(.A(G125), .B(G140), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n236), .B1(new_n558), .B2(new_n215), .ZN(new_n559));
  INV_X1    g373(.A(new_n237), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n542), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n544), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n238), .A2(KEYINPUT93), .A3(new_n542), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(new_n538), .B2(new_n539), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT19), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT19), .B1(new_n206), .B2(new_n209), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n215), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n217), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n526), .B2(new_n528), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n557), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n535), .ZN(new_n571));
  INV_X1    g385(.A(new_n528), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n217), .B(new_n567), .C1(new_n531), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n546), .A2(KEYINPUT94), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI211_X1 g389(.A(KEYINPUT20), .B(new_n556), .C1(new_n575), .C2(new_n547), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n571), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT94), .B1(new_n546), .B2(new_n573), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n547), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n577), .B1(new_n580), .B2(new_n555), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n554), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n248), .A2(G952), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n263), .B2(new_n353), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(G902), .B(G953), .C1(new_n263), .C2(new_n353), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(KEYINPUT98), .Z(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G217), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n393), .A2(new_n592), .A3(G953), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n305), .B2(G128), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n189), .A2(KEYINPUT97), .A3(G143), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT13), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G134), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n305), .A2(G128), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(G134), .A3(new_n600), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT96), .B1(new_n282), .B2(G122), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n608));
  INV_X1    g422(.A(G122), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(G116), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(G116), .B2(new_n609), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n612), .A2(G107), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(G107), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n604), .A2(new_n606), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n605), .A2(G134), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(KEYINPUT14), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(G107), .A3(new_n617), .ZN(new_n618));
  OAI221_X1 g432(.A(new_n611), .B1(KEYINPUT14), .B2(new_n400), .C1(G116), .C2(new_n609), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n603), .A2(new_n290), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n594), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n613), .A2(new_n614), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n606), .A2(new_n604), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n621), .A3(new_n593), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(G478), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT15), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n628), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n583), .A2(new_n591), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n521), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n277), .A2(new_n392), .A3(new_n462), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  NOR2_X1   g451(.A1(new_n266), .A2(new_n269), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n386), .A2(new_n455), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n639), .A2(G472), .B1(new_n389), .B2(new_n386), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n638), .A2(new_n275), .A3(new_n462), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n505), .A2(new_n514), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n519), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n623), .A2(new_n627), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT33), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n623), .A2(new_n647), .A3(new_n627), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(G478), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n629), .A2(new_n455), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n628), .B2(new_n629), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n582), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n644), .A2(new_n653), .A3(new_n590), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n642), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT99), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  NAND2_X1  g472(.A1(new_n632), .A2(new_n554), .ZN(new_n659));
  INV_X1    g473(.A(new_n581), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n580), .A2(new_n577), .A3(new_n555), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(KEYINPUT100), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n576), .B2(new_n581), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n659), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n519), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n505), .B2(new_n514), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n665), .A2(new_n591), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n642), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NAND2_X1  g485(.A1(new_n267), .A2(KEYINPUT25), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n259), .A3(new_n273), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n262), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n268), .A2(KEYINPUT83), .A3(new_n259), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n244), .A2(new_n246), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n251), .A2(KEYINPUT36), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT101), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n274), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n635), .A3(new_n462), .A4(new_n640), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n586), .B1(new_n588), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(new_n665), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n456), .A2(new_n461), .ZN(new_n691));
  INV_X1    g505(.A(new_n395), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n691), .A2(new_n692), .A3(new_n667), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n690), .A2(new_n693), .A3(new_n392), .A4(new_n681), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  XOR2_X1   g509(.A(new_n686), .B(KEYINPUT39), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n462), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n515), .A2(new_n518), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT38), .Z(new_n701));
  NOR3_X1   g515(.A1(new_n365), .A2(new_n366), .A3(new_n358), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n370), .A2(new_n369), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n455), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n390), .B2(new_n391), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n583), .A2(new_n633), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(KEYINPUT103), .A3(new_n519), .A4(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n519), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n711), .B1(new_n681), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n699), .A2(new_n707), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NAND3_X1  g529(.A1(new_n582), .A2(new_n652), .A3(new_n687), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n693), .A2(new_n392), .A3(new_n681), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND2_X1  g534(.A1(KEYINPUT105), .A2(G469), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n453), .A2(new_n455), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n453), .B2(new_n455), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n395), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n277), .A2(new_n724), .A3(new_n392), .A4(new_n654), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NAND4_X1  g541(.A1(new_n277), .A2(new_n724), .A3(new_n392), .A4(new_n668), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  INV_X1    g543(.A(new_n634), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n392), .A2(new_n681), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n722), .A2(new_n723), .A3(new_n644), .A4(new_n395), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND3_X1  g549(.A1(new_n674), .A2(new_n275), .A3(new_n675), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n377), .B1(new_n383), .B2(new_n385), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n389), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n378), .A2(new_n380), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n382), .A2(new_n357), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n384), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n702), .A2(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(G902), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT106), .B(G472), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n738), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT107), .B1(new_n736), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n639), .A2(new_n745), .B1(new_n389), .B2(new_n737), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n638), .A2(new_n749), .A3(new_n275), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n644), .A2(new_n583), .A3(new_n590), .A4(new_n633), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n724), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n752), .A2(KEYINPUT108), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT109), .B(G122), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G24));
  NAND4_X1  g576(.A1(new_n733), .A2(new_n681), .A3(new_n718), .A4(new_n750), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  NAND2_X1  g578(.A1(new_n386), .A2(new_n389), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT32), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(new_n767), .B1(G472), .B2(new_n374), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n736), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n666), .B1(new_n515), .B2(new_n518), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n691), .A2(new_n692), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n718), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n768), .A2(new_n771), .A3(new_n736), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n718), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NAND2_X1  g593(.A1(new_n277), .A2(new_n392), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n662), .A2(new_n664), .ZN(new_n781));
  INV_X1    g595(.A(new_n659), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n687), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT102), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n687), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n780), .A2(new_n787), .A3(new_n771), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n290), .ZN(G36));
  OAI21_X1  g603(.A(G469), .B1(new_n460), .B2(KEYINPUT45), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n459), .A2(new_n429), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n449), .A2(new_n442), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n460), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n790), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n457), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n456), .B1(new_n799), .B2(KEYINPUT46), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n798), .A2(new_n801), .A3(new_n457), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n692), .B(new_n696), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n770), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n583), .A2(new_n652), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n583), .A2(KEYINPUT43), .A3(new_n652), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n813), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT113), .A3(new_n811), .A4(new_n810), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n708), .A2(new_n640), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT44), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n814), .A2(new_n816), .A3(new_n817), .A4(KEYINPUT44), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n805), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G137), .ZN(G39));
  XNOR2_X1  g637(.A(new_n716), .B(KEYINPUT104), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n277), .A2(new_n824), .A3(new_n392), .A4(new_n804), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n692), .B1(new_n800), .B2(new_n802), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT47), .B(new_n692), .C1(new_n800), .C2(new_n802), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n825), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  NOR2_X1   g646(.A1(new_n722), .A2(new_n723), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n701), .B1(new_n834), .B2(KEYINPUT49), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n692), .A2(new_n520), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n706), .A2(new_n736), .A3(new_n807), .A4(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n835), .B(new_n837), .C1(KEYINPUT49), .C2(new_n834), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n828), .A2(new_n830), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n692), .B2(new_n834), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n815), .A2(new_n811), .A3(new_n810), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n586), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n752), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n804), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n701), .A2(new_n519), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n847), .A3(new_n724), .A4(new_n752), .ZN(new_n848));
  NOR2_X1   g662(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n724), .A2(new_n770), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n708), .A2(new_n747), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n853), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n851), .A2(new_n736), .A3(new_n585), .A4(new_n706), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n582), .A2(new_n652), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n846), .A2(new_n850), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n846), .A2(KEYINPUT51), .A3(new_n850), .A4(new_n861), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n842), .A2(new_n780), .A3(new_n851), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n858), .A2(new_n582), .A3(new_n652), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n584), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n724), .A2(new_n667), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n844), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n864), .A2(new_n865), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n725), .A2(new_n728), .A3(new_n682), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n515), .A2(new_n518), .A3(new_n520), .A4(new_n591), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT114), .B1(new_n582), .B2(new_n652), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n582), .A2(KEYINPUT114), .A3(new_n652), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n277), .A2(new_n880), .A3(new_n462), .A4(new_n640), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n636), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n583), .A2(new_n632), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n870), .A2(new_n731), .B1(new_n641), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n881), .A2(new_n636), .A3(KEYINPUT115), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n876), .A2(new_n884), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n392), .A2(new_n681), .A3(new_n785), .A4(new_n786), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n718), .A2(new_n392), .A3(new_n681), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n693), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n644), .A2(new_n583), .A3(new_n633), .A4(new_n686), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n708), .A2(new_n462), .A3(new_n706), .A4(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(KEYINPUT52), .A3(new_n763), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n694), .A2(new_n763), .A3(new_n719), .A4(new_n897), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n633), .A2(new_n554), .A3(new_n687), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n392), .A2(new_n681), .A3(new_n781), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n718), .A2(new_n681), .A3(new_n750), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n771), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n788), .B(new_n906), .C1(new_n775), .C2(new_n777), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n892), .A2(new_n902), .A3(new_n907), .A4(new_n760), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n906), .ZN(new_n911));
  INV_X1    g725(.A(new_n788), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT42), .B1(new_n776), .B2(new_n718), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n780), .A2(new_n774), .A3(new_n824), .A4(new_n771), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n911), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n757), .B(new_n754), .C1(new_n751), .C2(new_n748), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT108), .B1(new_n752), .B2(new_n755), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n891), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n920));
  NOR2_X1   g734(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n895), .A2(new_n763), .A3(new_n897), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n899), .A2(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT54), .B1(new_n910), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n908), .A2(new_n909), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n919), .A2(KEYINPUT53), .A3(new_n926), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(KEYINPUT117), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(KEYINPUT54), .C1(new_n910), .C2(new_n927), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n874), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(G952), .A2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n838), .B1(new_n936), .B2(new_n937), .ZN(G75));
  NAND2_X1  g752(.A1(new_n929), .A2(new_n930), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(G210), .A3(G902), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT56), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n511), .A2(new_n512), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT120), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n473), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n940), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n940), .B2(new_n941), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n248), .A2(G952), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(G51));
  XNOR2_X1  g763(.A(new_n457), .B(KEYINPUT57), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n931), .B1(new_n929), .B2(new_n930), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n453), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n939), .A2(G902), .A3(new_n798), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(G54));
  AND2_X1   g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT53), .B1(new_n919), .B2(new_n902), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT115), .B1(new_n881), .B2(new_n636), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n959), .A2(new_n875), .A3(new_n888), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n760), .A2(new_n960), .A3(new_n890), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n961), .A2(new_n925), .A3(new_n909), .A4(new_n915), .ZN(new_n962));
  OAI211_X1 g776(.A(G902), .B(new_n957), .C1(new_n958), .C2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n580), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n948), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n939), .A2(G902), .A3(new_n580), .A4(new_n957), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n965), .A2(KEYINPUT121), .A3(new_n966), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(G60));
  AND2_X1   g786(.A1(new_n646), .A2(new_n648), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n650), .B(KEYINPUT59), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n951), .B2(new_n952), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n966), .ZN(new_n977));
  INV_X1    g791(.A(new_n974), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n933), .A2(new_n935), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n973), .B2(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT60), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n939), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n272), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n948), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n929), .B2(new_n930), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n679), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n986), .B(new_n988), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n989));
  OAI211_X1 g803(.A(KEYINPUT122), .B(new_n966), .C1(new_n987), .C2(new_n272), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n966), .B1(new_n987), .B2(new_n272), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n939), .A2(new_n679), .A3(new_n983), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n990), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n994), .ZN(G66));
  OAI21_X1  g809(.A(G953), .B1(new_n589), .B2(new_n468), .ZN(new_n996));
  INV_X1    g810(.A(new_n961), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(G953), .ZN(new_n998));
  INV_X1    g812(.A(new_n943), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(G898), .B2(new_n248), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(G69));
  NAND3_X1  g815(.A1(new_n769), .A2(new_n667), .A3(new_n709), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n803), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT126), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1005), .B1(new_n803), .B2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n788), .B1(new_n775), .B2(new_n777), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1007), .A2(new_n831), .A3(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n694), .A2(new_n719), .A3(new_n763), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT125), .B1(new_n822), .B2(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n822), .A2(KEYINPUT125), .A3(new_n1010), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1009), .B(new_n248), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n565), .A2(new_n566), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT123), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n381), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n248), .B1(G227), .B2(G900), .ZN(new_n1019));
  AOI22_X1  g833(.A1(new_n1013), .A2(new_n1018), .B1(KEYINPUT127), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1019), .A2(KEYINPUT127), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n879), .A2(new_n878), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n804), .B1(new_n1022), .B2(new_n885), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n769), .A2(new_n1023), .A3(new_n462), .A4(new_n696), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n831), .A2(new_n822), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n714), .A2(new_n1010), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT62), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n714), .A2(new_n1010), .A3(KEYINPUT62), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(KEYINPUT124), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT124), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1025), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(G953), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1020), .B(new_n1021), .C1(new_n1035), .C2(new_n1016), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1034), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1033), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n248), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n1017), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1021), .B1(new_n1041), .B2(new_n1020), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1037), .A2(new_n1042), .ZN(G72));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  OAI21_X1  g859(.A(new_n1009), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1045), .B1(new_n1046), .B2(new_n961), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1047), .A2(new_n382), .A3(new_n358), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n910), .A2(new_n927), .ZN(new_n1049));
  INV_X1    g863(.A(new_n367), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1045), .B1(new_n1050), .B2(new_n702), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n1048), .B(new_n966), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1032), .A2(new_n997), .A3(new_n1034), .ZN(new_n1053));
  AOI211_X1 g867(.A(new_n382), .B(new_n358), .C1(new_n1053), .C2(new_n1045), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1052), .A2(new_n1054), .ZN(G57));
endmodule


