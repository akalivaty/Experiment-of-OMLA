

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764;

  XNOR2_X1 U369 ( .A(n640), .B(n466), .ZN(n679) );
  XNOR2_X1 U370 ( .A(n489), .B(G110), .ZN(n488) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n548) );
  XNOR2_X1 U372 ( .A(n737), .B(n413), .ZN(n546) );
  INV_X2 U373 ( .A(G953), .ZN(n748) );
  OR2_X1 U374 ( .A1(n486), .A2(n485), .ZN(n348) );
  XOR2_X1 U375 ( .A(n723), .B(n366), .Z(n349) );
  NOR2_X2 U376 ( .A1(n653), .A2(n729), .ZN(n656) );
  OR2_X2 U377 ( .A1(n595), .A2(n471), .ZN(n354) );
  NOR2_X1 U378 ( .A1(G902), .A2(n723), .ZN(n531) );
  NAND2_X1 U379 ( .A1(n439), .A2(n348), .ZN(n663) );
  NOR2_X1 U380 ( .A1(n568), .A2(n440), .ZN(n569) );
  INV_X1 U381 ( .A(n707), .ZN(n432) );
  INV_X1 U382 ( .A(n605), .ZN(n448) );
  NAND2_X2 U383 ( .A1(n622), .A2(n506), .ZN(n507) );
  INV_X1 U384 ( .A(KEYINPUT18), .ZN(n437) );
  INV_X1 U385 ( .A(KEYINPUT16), .ZN(n489) );
  AND2_X1 U386 ( .A1(n453), .A2(n354), .ZN(n480) );
  AND2_X1 U387 ( .A1(n395), .A2(n394), .ZN(n388) );
  AND2_X1 U388 ( .A1(n468), .A2(n444), .ZN(n453) );
  AND2_X1 U389 ( .A1(n399), .A2(n359), .ZN(n397) );
  XNOR2_X1 U390 ( .A(KEYINPUT114), .B(n633), .ZN(n757) );
  NOR2_X1 U391 ( .A1(n545), .A2(n567), .ZN(n570) );
  OR2_X1 U392 ( .A1(n683), .A2(n682), .ZN(n465) );
  AND2_X1 U393 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U394 ( .A(n547), .B(n472), .ZN(n720) );
  XNOR2_X1 U395 ( .A(n411), .B(n410), .ZN(n409) );
  NAND2_X1 U396 ( .A1(n512), .A2(n511), .ZN(n538) );
  XNOR2_X1 U397 ( .A(n501), .B(n356), .ZN(n411) );
  NAND2_X1 U398 ( .A1(n509), .A2(n508), .ZN(n512) );
  XNOR2_X1 U399 ( .A(n499), .B(n509), .ZN(n410) );
  XNOR2_X1 U400 ( .A(n437), .B(KEYINPUT17), .ZN(n436) );
  XNOR2_X1 U401 ( .A(G143), .B(G131), .ZN(n523) );
  INV_X1 U402 ( .A(G134), .ZN(n508) );
  XNOR2_X1 U403 ( .A(n416), .B(n363), .ZN(n653) );
  NOR2_X1 U404 ( .A1(n711), .A2(n365), .ZN(n416) );
  BUF_X1 U405 ( .A(n599), .Z(n640) );
  AND2_X2 U406 ( .A1(n575), .A2(n688), .ZN(n584) );
  BUF_X1 U407 ( .A(n668), .Z(n350) );
  XNOR2_X1 U408 ( .A(G146), .B(G125), .ZN(n518) );
  NAND2_X1 U409 ( .A1(n351), .A2(n679), .ZN(n377) );
  OR2_X1 U410 ( .A1(n441), .A2(n613), .ZN(n376) );
  NAND2_X2 U411 ( .A1(n405), .A2(n402), .ZN(n616) );
  NAND2_X1 U412 ( .A1(n544), .A2(n404), .ZN(n403) );
  INV_X1 U413 ( .A(G475), .ZN(n430) );
  INV_X1 U414 ( .A(G210), .ZN(n431) );
  INV_X1 U415 ( .A(KEYINPUT83), .ZN(n471) );
  NAND2_X1 U416 ( .A1(n748), .A2(G224), .ZN(n447) );
  XNOR2_X1 U417 ( .A(n460), .B(n362), .ZN(n395) );
  NAND2_X1 U418 ( .A1(n423), .A2(n663), .ZN(n435) );
  NAND2_X1 U419 ( .A1(n720), .A2(G469), .ZN(n407) );
  XNOR2_X1 U420 ( .A(n566), .B(n565), .ZN(n690) );
  XOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n550) );
  XNOR2_X1 U422 ( .A(n523), .B(n522), .ZN(n524) );
  INV_X1 U423 ( .A(KEYINPUT99), .ZN(n522) );
  XNOR2_X1 U424 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n519) );
  OR2_X1 U425 ( .A1(G237), .A2(G902), .ZN(n504) );
  NAND2_X1 U426 ( .A1(n377), .A2(n378), .ZN(n375) );
  INV_X1 U427 ( .A(n377), .ZN(n373) );
  NOR2_X1 U428 ( .A1(n585), .A2(KEYINPUT34), .ZN(n400) );
  AND2_X1 U429 ( .A1(n458), .A2(n612), .ZN(n441) );
  NOR2_X1 U430 ( .A1(n545), .A2(n485), .ZN(n482) );
  NAND2_X1 U431 ( .A1(n545), .A2(n485), .ZN(n484) );
  OR2_X1 U432 ( .A1(n652), .A2(G902), .ZN(n450) );
  XNOR2_X1 U433 ( .A(n383), .B(n433), .ZN(n561) );
  INV_X1 U434 ( .A(KEYINPUT8), .ZN(n433) );
  XNOR2_X1 U435 ( .A(n543), .B(n542), .ZN(n474) );
  INV_X1 U436 ( .A(G107), .ZN(n542) );
  XNOR2_X1 U437 ( .A(G110), .B(G104), .ZN(n543) );
  XOR2_X1 U438 ( .A(KEYINPUT67), .B(G101), .Z(n539) );
  XOR2_X1 U439 ( .A(G137), .B(G140), .Z(n556) );
  XNOR2_X1 U440 ( .A(n457), .B(n456), .ZN(n624) );
  INV_X1 U441 ( .A(KEYINPUT110), .ZN(n456) );
  OR2_X1 U442 ( .A1(n618), .A2(n617), .ZN(n457) );
  XNOR2_X1 U443 ( .A(n434), .B(G478), .ZN(n591) );
  NOR2_X1 U444 ( .A1(n725), .A2(G902), .ZN(n434) );
  INV_X1 U445 ( .A(KEYINPUT104), .ZN(n485) );
  INV_X1 U446 ( .A(KEYINPUT2), .ZN(n370) );
  NOR2_X1 U447 ( .A1(n471), .A2(KEYINPUT44), .ZN(n469) );
  AND2_X1 U448 ( .A1(n471), .A2(KEYINPUT44), .ZN(n470) );
  INV_X1 U449 ( .A(KEYINPUT38), .ZN(n466) );
  INV_X1 U450 ( .A(G902), .ZN(n404) );
  NAND2_X1 U451 ( .A1(G469), .A2(G902), .ZN(n406) );
  XNOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n500) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n491) );
  NAND2_X1 U454 ( .A1(n385), .A2(KEYINPUT48), .ZN(n384) );
  INV_X1 U455 ( .A(KEYINPUT65), .ZN(n479) );
  INV_X1 U456 ( .A(KEYINPUT82), .ZN(n477) );
  INV_X1 U457 ( .A(KEYINPUT28), .ZN(n442) );
  NAND2_X1 U458 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U459 ( .A1(n588), .A2(n590), .ZN(n532) );
  NAND2_X1 U460 ( .A1(n448), .A2(n355), .ZN(n628) );
  NOR2_X1 U461 ( .A1(n682), .A2(n691), .ZN(n536) );
  XOR2_X1 U462 ( .A(n610), .B(n451), .Z(n351) );
  XNOR2_X1 U463 ( .A(n452), .B(KEYINPUT30), .ZN(n451) );
  INV_X1 U464 ( .A(KEYINPUT107), .ZN(n452) );
  NOR2_X1 U465 ( .A1(n691), .A2(n690), .ZN(n688) );
  INV_X1 U466 ( .A(G472), .ZN(n429) );
  XNOR2_X1 U467 ( .A(n555), .B(n554), .ZN(n652) );
  XNOR2_X1 U468 ( .A(n547), .B(n546), .ZN(n555) );
  XNOR2_X1 U469 ( .A(G137), .B(G113), .ZN(n552) );
  XNOR2_X1 U470 ( .A(n559), .B(n381), .ZN(n380) );
  XNOR2_X1 U471 ( .A(KEYINPUT93), .B(KEYINPUT24), .ZN(n559) );
  XNOR2_X1 U472 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n381) );
  XNOR2_X1 U473 ( .A(G128), .B(G119), .ZN(n558) );
  XNOR2_X1 U474 ( .A(n529), .B(n528), .ZN(n723) );
  XNOR2_X1 U475 ( .A(G902), .B(KEYINPUT15), .ZN(n650) );
  NAND2_X1 U476 ( .A1(n357), .A2(n372), .ZN(n648) );
  NAND2_X1 U477 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U478 ( .A1(n441), .A2(n351), .ZN(n641) );
  NOR2_X1 U479 ( .A1(n482), .A2(n694), .ZN(n481) );
  XNOR2_X1 U480 ( .A(n580), .B(KEYINPUT96), .ZN(n611) );
  AND2_X1 U481 ( .A1(n616), .A2(n688), .ZN(n580) );
  INV_X1 U482 ( .A(KEYINPUT0), .ZN(n475) );
  INV_X1 U483 ( .A(KEYINPUT3), .ZN(n463) );
  XNOR2_X1 U484 ( .A(n459), .B(n742), .ZN(n728) );
  XNOR2_X1 U485 ( .A(n382), .B(n379), .ZN(n459) );
  NAND2_X1 U486 ( .A1(n561), .A2(G221), .ZN(n382) );
  XNOR2_X1 U487 ( .A(n560), .B(n380), .ZN(n379) );
  XOR2_X1 U488 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n515) );
  XNOR2_X1 U489 ( .A(n541), .B(n473), .ZN(n472) );
  XNOR2_X1 U490 ( .A(n474), .B(n540), .ZN(n473) );
  XNOR2_X1 U491 ( .A(n614), .B(KEYINPUT40), .ZN(n761) );
  NAND2_X1 U492 ( .A1(n648), .A2(n350), .ZN(n614) );
  INV_X1 U493 ( .A(KEYINPUT60), .ZN(n417) );
  INV_X1 U494 ( .A(KEYINPUT56), .ZN(n419) );
  XNOR2_X1 U495 ( .A(n667), .B(n467), .ZN(G30) );
  INV_X1 U496 ( .A(G128), .ZN(n467) );
  OR2_X1 U497 ( .A1(n657), .A2(n469), .ZN(n352) );
  XNOR2_X1 U498 ( .A(n592), .B(KEYINPUT101), .ZN(n668) );
  XOR2_X1 U499 ( .A(KEYINPUT4), .B(G131), .Z(n353) );
  XNOR2_X1 U500 ( .A(n518), .B(n519), .ZN(n557) );
  AND2_X1 U501 ( .A1(n615), .A2(n350), .ZN(n355) );
  XOR2_X1 U502 ( .A(n447), .B(n498), .Z(n356) );
  BUF_X1 U503 ( .A(n609), .Z(n694) );
  INV_X1 U504 ( .A(n690), .ZN(n440) );
  AND2_X1 U505 ( .A1(n376), .A2(n375), .ZN(n357) );
  AND2_X1 U506 ( .A1(n593), .A2(n625), .ZN(n358) );
  AND2_X1 U507 ( .A1(n398), .A2(n578), .ZN(n359) );
  AND2_X1 U508 ( .A1(n481), .A2(n690), .ZN(n360) );
  XOR2_X1 U509 ( .A(n537), .B(KEYINPUT66), .Z(n361) );
  INV_X1 U510 ( .A(n613), .ZN(n378) );
  XNOR2_X1 U511 ( .A(KEYINPUT81), .B(KEYINPUT39), .ZN(n613) );
  INV_X1 U512 ( .A(n729), .ZN(n424) );
  XOR2_X1 U513 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n362) );
  XOR2_X1 U514 ( .A(n652), .B(n651), .Z(n363) );
  XNOR2_X1 U515 ( .A(n718), .B(n717), .ZN(n364) );
  INV_X1 U516 ( .A(KEYINPUT48), .ZN(n394) );
  OR2_X1 U517 ( .A1(n650), .A2(n429), .ZN(n365) );
  XNOR2_X1 U518 ( .A(KEYINPUT59), .B(KEYINPUT87), .ZN(n366) );
  OR2_X1 U519 ( .A1(n650), .A2(n430), .ZN(n367) );
  OR2_X1 U520 ( .A1(n650), .A2(n431), .ZN(n368) );
  XNOR2_X1 U521 ( .A(n727), .B(n728), .ZN(n414) );
  NAND2_X1 U522 ( .A1(n428), .A2(n427), .ZN(n371) );
  XNOR2_X1 U523 ( .A(n598), .B(KEYINPUT45), .ZN(n428) );
  NOR2_X1 U524 ( .A1(n369), .A2(n729), .ZN(G54) );
  XNOR2_X1 U525 ( .A(n722), .B(n721), .ZN(n369) );
  XNOR2_X2 U526 ( .A(n371), .B(n370), .ZN(n711) );
  AND2_X1 U527 ( .A1(n441), .A2(n613), .ZN(n374) );
  NAND2_X1 U528 ( .A1(n748), .A2(G234), .ZN(n383) );
  NAND2_X1 U529 ( .A1(n386), .A2(n384), .ZN(n392) );
  INV_X1 U530 ( .A(n387), .ZN(n385) );
  NAND2_X1 U531 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U532 ( .A(n462), .B(n461), .ZN(n387) );
  NOR2_X1 U533 ( .A1(n392), .A2(n389), .ZN(n649) );
  NAND2_X1 U534 ( .A1(n390), .A2(n393), .ZN(n389) );
  NAND2_X1 U535 ( .A1(n391), .A2(KEYINPUT48), .ZN(n390) );
  INV_X1 U536 ( .A(n395), .ZN(n391) );
  INV_X1 U537 ( .A(n677), .ZN(n393) );
  NAND2_X1 U538 ( .A1(n397), .A2(n396), .ZN(n579) );
  NAND2_X1 U539 ( .A1(n708), .A2(KEYINPUT34), .ZN(n396) );
  NAND2_X1 U540 ( .A1(n585), .A2(KEYINPUT34), .ZN(n398) );
  NAND2_X1 U541 ( .A1(n401), .A2(n400), .ZN(n399) );
  INV_X1 U542 ( .A(n708), .ZN(n401) );
  XNOR2_X2 U543 ( .A(n577), .B(KEYINPUT33), .ZN(n708) );
  XNOR2_X2 U544 ( .A(n616), .B(KEYINPUT1), .ZN(n575) );
  OR2_X1 U545 ( .A1(n720), .A2(n403), .ZN(n402) );
  XNOR2_X2 U546 ( .A(n408), .B(n527), .ZN(n735) );
  XNOR2_X2 U547 ( .A(n513), .B(n488), .ZN(n408) );
  XNOR2_X2 U548 ( .A(n412), .B(n409), .ZN(n718) );
  XNOR2_X2 U549 ( .A(n735), .B(n546), .ZN(n412) );
  INV_X1 U550 ( .A(n539), .ZN(n413) );
  XNOR2_X2 U551 ( .A(n464), .B(n463), .ZN(n737) );
  XNOR2_X2 U552 ( .A(n487), .B(G122), .ZN(n527) );
  NOR2_X1 U553 ( .A1(n414), .A2(n729), .ZN(G66) );
  XNOR2_X1 U554 ( .A(n426), .B(n349), .ZN(n425) );
  OR2_X2 U555 ( .A1(n711), .A2(n368), .ZN(n422) );
  NOR2_X1 U556 ( .A1(n415), .A2(n729), .ZN(G63) );
  XNOR2_X1 U557 ( .A(n724), .B(n725), .ZN(n415) );
  XNOR2_X1 U558 ( .A(n418), .B(n417), .ZN(G60) );
  NAND2_X1 U559 ( .A1(n425), .A2(n424), .ZN(n418) );
  XNOR2_X1 U560 ( .A(n420), .B(n419), .ZN(G51) );
  NAND2_X1 U561 ( .A1(n421), .A2(n424), .ZN(n420) );
  XNOR2_X1 U562 ( .A(n422), .B(n364), .ZN(n421) );
  XNOR2_X1 U563 ( .A(n423), .B(G119), .ZN(G21) );
  XNOR2_X2 U564 ( .A(n571), .B(KEYINPUT32), .ZN(n423) );
  OR2_X2 U565 ( .A1(n711), .A2(n367), .ZN(n426) );
  INV_X1 U566 ( .A(n747), .ZN(n427) );
  AND2_X1 U567 ( .A1(n428), .A2(n748), .ZN(n733) );
  NOR2_X1 U568 ( .A1(n711), .A2(n650), .ZN(n726) );
  NAND2_X1 U569 ( .A1(n432), .A2(n624), .ZN(n620) );
  XNOR2_X2 U570 ( .A(n465), .B(n619), .ZN(n707) );
  XNOR2_X1 U571 ( .A(n517), .B(n538), .ZN(n445) );
  NAND2_X1 U572 ( .A1(n761), .A2(n763), .ZN(n460) );
  XNOR2_X2 U573 ( .A(n435), .B(KEYINPUT84), .ZN(n594) );
  NOR2_X2 U574 ( .A1(n605), .A2(n576), .ZN(n577) );
  XNOR2_X1 U575 ( .A(n500), .B(n436), .ZN(n501) );
  INV_X1 U576 ( .A(n438), .ZN(n439) );
  NAND2_X1 U577 ( .A1(n483), .A2(n360), .ZN(n438) );
  INV_X1 U578 ( .A(n518), .ZN(n499) );
  NAND2_X1 U579 ( .A1(n581), .A2(n536), .ZN(n446) );
  XNOR2_X2 U580 ( .A(n507), .B(n475), .ZN(n581) );
  NAND2_X1 U581 ( .A1(n690), .A2(n612), .ZN(n604) );
  XNOR2_X1 U582 ( .A(n443), .B(n442), .ZN(n618) );
  AND2_X1 U583 ( .A1(n615), .A2(n609), .ZN(n443) );
  XNOR2_X1 U584 ( .A(n611), .B(KEYINPUT106), .ZN(n458) );
  NOR2_X1 U585 ( .A1(n352), .A2(n358), .ZN(n444) );
  NAND2_X1 U586 ( .A1(n594), .A2(KEYINPUT44), .ZN(n572) );
  XNOR2_X1 U587 ( .A(n445), .B(n516), .ZN(n725) );
  INV_X2 U588 ( .A(G116), .ZN(n490) );
  OR2_X2 U589 ( .A1(n568), .A2(n484), .ZN(n483) );
  XNOR2_X2 U590 ( .A(n446), .B(n361), .ZN(n568) );
  INV_X2 U591 ( .A(n510), .ZN(n509) );
  INV_X1 U592 ( .A(n628), .ZN(n626) );
  XNOR2_X1 U593 ( .A(n557), .B(n449), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(n449) );
  XNOR2_X2 U595 ( .A(n627), .B(n505), .ZN(n622) );
  NAND2_X2 U596 ( .A1(n599), .A2(n678), .ZN(n627) );
  XNOR2_X2 U597 ( .A(n450), .B(G472), .ZN(n609) );
  XNOR2_X1 U598 ( .A(n454), .B(n477), .ZN(n476) );
  NAND2_X1 U599 ( .A1(n478), .A2(n480), .ZN(n454) );
  NAND2_X1 U600 ( .A1(n455), .A2(KEYINPUT47), .ZN(n634) );
  NAND2_X1 U601 ( .A1(n669), .A2(n625), .ZN(n455) );
  XNOR2_X1 U602 ( .A(n513), .B(G122), .ZN(n514) );
  XNOR2_X2 U603 ( .A(n490), .B(G107), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n572), .B(n479), .ZN(n478) );
  NAND2_X1 U605 ( .A1(n476), .A2(n597), .ZN(n598) );
  NOR2_X1 U606 ( .A1(n728), .A2(G902), .ZN(n566) );
  INV_X1 U607 ( .A(KEYINPUT69), .ZN(n461) );
  AND2_X1 U608 ( .A1(n646), .A2(n762), .ZN(n462) );
  XNOR2_X2 U609 ( .A(KEYINPUT70), .B(G119), .ZN(n464) );
  NAND2_X1 U610 ( .A1(n595), .A2(n470), .ZN(n468) );
  XNOR2_X2 U611 ( .A(n579), .B(KEYINPUT35), .ZN(n595) );
  XNOR2_X2 U612 ( .A(n744), .B(G146), .ZN(n547) );
  XNOR2_X2 U613 ( .A(n538), .B(n353), .ZN(n744) );
  NAND2_X1 U614 ( .A1(n486), .A2(n545), .ZN(n574) );
  INV_X1 U615 ( .A(n568), .ZN(n486) );
  XNOR2_X2 U616 ( .A(G113), .B(G104), .ZN(n487) );
  XNOR2_X2 U617 ( .A(G143), .B(G128), .ZN(n510) );
  XNOR2_X2 U618 ( .A(n609), .B(KEYINPUT6), .ZN(n605) );
  INV_X1 U619 ( .A(KEYINPUT77), .ZN(n498) );
  XNOR2_X1 U620 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U621 ( .A(n654), .B(KEYINPUT88), .ZN(n655) );
  NOR2_X1 U622 ( .A1(G952), .A2(n748), .ZN(n729) );
  XNOR2_X1 U623 ( .A(n491), .B(KEYINPUT14), .ZN(n492) );
  XNOR2_X1 U624 ( .A(KEYINPUT74), .B(n492), .ZN(n495) );
  NAND2_X1 U625 ( .A1(n495), .A2(G902), .ZN(n493) );
  XOR2_X1 U626 ( .A(KEYINPUT91), .B(n493), .Z(n600) );
  INV_X1 U627 ( .A(n600), .ZN(n494) );
  NOR2_X1 U628 ( .A1(G898), .A2(n748), .ZN(n739) );
  NAND2_X1 U629 ( .A1(n494), .A2(n739), .ZN(n497) );
  NAND2_X1 U630 ( .A1(G952), .A2(n495), .ZN(n706) );
  NOR2_X1 U631 ( .A1(G953), .A2(n706), .ZN(n496) );
  XOR2_X1 U632 ( .A(KEYINPUT90), .B(n496), .Z(n603) );
  NAND2_X1 U633 ( .A1(n497), .A2(n603), .ZN(n506) );
  NAND2_X1 U634 ( .A1(n718), .A2(n650), .ZN(n503) );
  AND2_X1 U635 ( .A1(G210), .A2(n504), .ZN(n502) );
  XNOR2_X2 U636 ( .A(n503), .B(n502), .ZN(n599) );
  NAND2_X1 U637 ( .A1(G214), .A2(n504), .ZN(n678) );
  XNOR2_X1 U638 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n505) );
  NAND2_X1 U639 ( .A1(G134), .A2(n510), .ZN(n511) );
  NAND2_X1 U640 ( .A1(n561), .A2(G217), .ZN(n517) );
  XNOR2_X1 U641 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U642 ( .A(n591), .ZN(n588) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n521) );
  XNOR2_X1 U644 ( .A(G140), .B(KEYINPUT100), .ZN(n520) );
  XNOR2_X1 U645 ( .A(n521), .B(n520), .ZN(n525) );
  NAND2_X1 U646 ( .A1(G214), .A2(n548), .ZN(n526) );
  XNOR2_X1 U647 ( .A(KEYINPUT13), .B(G475), .ZN(n530) );
  XNOR2_X1 U648 ( .A(n531), .B(n530), .ZN(n590) );
  XNOR2_X1 U649 ( .A(n532), .B(KEYINPUT103), .ZN(n682) );
  XOR2_X1 U650 ( .A(KEYINPUT21), .B(KEYINPUT95), .Z(n535) );
  NAND2_X1 U651 ( .A1(G234), .A2(n650), .ZN(n533) );
  XNOR2_X1 U652 ( .A(KEYINPUT20), .B(n533), .ZN(n562) );
  NAND2_X1 U653 ( .A1(n562), .A2(G221), .ZN(n534) );
  XNOR2_X1 U654 ( .A(n535), .B(n534), .ZN(n691) );
  XNOR2_X1 U655 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n537) );
  XNOR2_X1 U656 ( .A(n539), .B(n556), .ZN(n541) );
  NAND2_X1 U657 ( .A1(G227), .A2(n748), .ZN(n540) );
  INV_X1 U658 ( .A(G469), .ZN(n544) );
  INV_X1 U659 ( .A(n575), .ZN(n545) );
  NAND2_X1 U660 ( .A1(n548), .A2(G210), .ZN(n549) );
  XNOR2_X1 U661 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U662 ( .A(n551), .B(G116), .Z(n553) );
  XNOR2_X1 U663 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U664 ( .A(n557), .B(n556), .ZN(n742) );
  XNOR2_X1 U665 ( .A(n558), .B(G110), .ZN(n560) );
  XOR2_X1 U666 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n564) );
  NAND2_X1 U667 ( .A1(G217), .A2(n562), .ZN(n563) );
  XNOR2_X1 U668 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U669 ( .A(KEYINPUT79), .B(n605), .ZN(n567) );
  NAND2_X1 U670 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U671 ( .A1(n440), .A2(n605), .ZN(n573) );
  NOR2_X1 U672 ( .A1(n574), .A2(n573), .ZN(n657) );
  XNOR2_X1 U673 ( .A(n584), .B(KEYINPUT105), .ZN(n576) );
  INV_X1 U674 ( .A(n581), .ZN(n585) );
  INV_X1 U675 ( .A(n590), .ZN(n589) );
  NOR2_X1 U676 ( .A1(n589), .A2(n591), .ZN(n644) );
  XNOR2_X1 U677 ( .A(n644), .B(KEYINPUT78), .ZN(n578) );
  NAND2_X1 U678 ( .A1(n611), .A2(n581), .ZN(n582) );
  NOR2_X1 U679 ( .A1(n582), .A2(n694), .ZN(n583) );
  XNOR2_X1 U680 ( .A(n583), .B(KEYINPUT97), .ZN(n659) );
  NAND2_X1 U681 ( .A1(n694), .A2(n584), .ZN(n699) );
  NOR2_X1 U682 ( .A1(n585), .A2(n699), .ZN(n587) );
  XNOR2_X1 U683 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n586) );
  XNOR2_X1 U684 ( .A(n587), .B(n586), .ZN(n674) );
  NAND2_X1 U685 ( .A1(n659), .A2(n674), .ZN(n593) );
  NAND2_X1 U686 ( .A1(n589), .A2(n588), .ZN(n673) );
  XOR2_X1 U687 ( .A(KEYINPUT102), .B(n673), .Z(n647) );
  NAND2_X1 U688 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U689 ( .A1(n647), .A2(n350), .ZN(n684) );
  INV_X1 U690 ( .A(n684), .ZN(n625) );
  NOR2_X1 U691 ( .A1(n594), .A2(KEYINPUT44), .ZN(n596) );
  INV_X1 U692 ( .A(n595), .ZN(n760) );
  NAND2_X1 U693 ( .A1(n596), .A2(n760), .ZN(n597) );
  NOR2_X1 U694 ( .A1(G900), .A2(n600), .ZN(n601) );
  NAND2_X1 U695 ( .A1(G953), .A2(n601), .ZN(n602) );
  NAND2_X1 U696 ( .A1(n603), .A2(n602), .ZN(n612) );
  NOR2_X1 U697 ( .A1(n691), .A2(n604), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n626), .A2(n678), .ZN(n606) );
  NOR2_X1 U699 ( .A1(n575), .A2(n606), .ZN(n607) );
  XNOR2_X1 U700 ( .A(n607), .B(KEYINPUT43), .ZN(n608) );
  NOR2_X1 U701 ( .A1(n640), .A2(n608), .ZN(n677) );
  NAND2_X1 U702 ( .A1(n678), .A2(n609), .ZN(n610) );
  XNOR2_X1 U703 ( .A(n616), .B(KEYINPUT109), .ZN(n617) );
  XNOR2_X1 U704 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n619) );
  XNOR2_X1 U705 ( .A(n620), .B(KEYINPUT42), .ZN(n621) );
  XNOR2_X1 U706 ( .A(KEYINPUT112), .B(n621), .ZN(n763) );
  BUF_X1 U707 ( .A(n622), .Z(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n664) );
  INV_X1 U709 ( .A(n664), .ZN(n669) );
  NOR2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n631) );
  XNOR2_X1 U711 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT113), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n631), .B(n630), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n575), .A2(n632), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n757), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n684), .A2(KEYINPUT47), .ZN(n635) );
  XNOR2_X1 U717 ( .A(n635), .B(KEYINPUT73), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n664), .A2(n636), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n637), .B(KEYINPUT72), .ZN(n638) );
  NOR2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n646) );
  INV_X1 U721 ( .A(n640), .ZN(n642) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U724 ( .A(KEYINPUT108), .B(n645), .ZN(n762) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n676) );
  NAND2_X1 U726 ( .A1(n649), .A2(n676), .ZN(n747) );
  XOR2_X1 U727 ( .A(KEYINPUT62), .B(KEYINPUT115), .Z(n651) );
  XOR2_X1 U728 ( .A(KEYINPUT63), .B(KEYINPUT116), .Z(n654) );
  XNOR2_X1 U729 ( .A(n656), .B(n655), .ZN(G57) );
  XOR2_X1 U730 ( .A(G101), .B(n657), .Z(G3) );
  INV_X1 U731 ( .A(n350), .ZN(n671) );
  NOR2_X1 U732 ( .A1(n671), .A2(n659), .ZN(n658) );
  XOR2_X1 U733 ( .A(G104), .B(n658), .Z(G6) );
  NOR2_X1 U734 ( .A1(n673), .A2(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U737 ( .A(G107), .B(n662), .ZN(G9) );
  XNOR2_X1 U738 ( .A(n663), .B(G110), .ZN(G12) );
  XOR2_X1 U739 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n666) );
  OR2_X1 U740 ( .A1(n664), .A2(n673), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n669), .A2(n350), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n670), .B(G146), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n674), .A2(n671), .ZN(n672) );
  XOR2_X1 U745 ( .A(G113), .B(n672), .Z(G15) );
  NOR2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U747 ( .A(G116), .B(n675), .Z(G18) );
  XNOR2_X1 U748 ( .A(G134), .B(n676), .ZN(G36) );
  XOR2_X1 U749 ( .A(G140), .B(n677), .Z(G42) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT120), .ZN(n681) );
  NOR2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n687), .A2(n708), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n688), .A2(n575), .ZN(n689) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(n689), .Z(n697) );
  XOR2_X1 U758 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n693) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n693), .B(n692), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n707), .A2(n701), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n713), .A2(G953), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n714), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U774 ( .A(KEYINPUT86), .B(KEYINPUT80), .Z(n716) );
  XNOR2_X1 U775 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n715) );
  XNOR2_X1 U776 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U777 ( .A1(n726), .A2(G469), .ZN(n722) );
  XOR2_X1 U778 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  XNOR2_X1 U779 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U780 ( .A1(G478), .A2(n726), .ZN(n724) );
  NAND2_X1 U781 ( .A1(G217), .A2(n726), .ZN(n727) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U783 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U784 ( .A1(n731), .A2(G898), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n732), .B(KEYINPUT121), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n741) );
  XOR2_X1 U787 ( .A(n735), .B(G101), .Z(n736) );
  XNOR2_X1 U788 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U790 ( .A(n741), .B(n740), .Z(G69) );
  XOR2_X1 U791 ( .A(n742), .B(KEYINPUT122), .Z(n743) );
  XNOR2_X1 U792 ( .A(n744), .B(n743), .ZN(n750) );
  INV_X1 U793 ( .A(n750), .ZN(n745) );
  XNOR2_X1 U794 ( .A(KEYINPUT123), .B(n745), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n756) );
  XNOR2_X1 U797 ( .A(G227), .B(n750), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n751), .B(KEYINPUT124), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U800 ( .A1(G953), .A2(n753), .ZN(n754) );
  XOR2_X1 U801 ( .A(KEYINPUT125), .B(n754), .Z(n755) );
  NAND2_X1 U802 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U803 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n759) );
  XNOR2_X1 U804 ( .A(n757), .B(G125), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n759), .B(n758), .ZN(G27) );
  XNOR2_X1 U806 ( .A(G122), .B(n760), .ZN(G24) );
  XNOR2_X1 U807 ( .A(n761), .B(G131), .ZN(G33) );
  XNOR2_X1 U808 ( .A(G143), .B(n762), .ZN(G45) );
  XNOR2_X1 U809 ( .A(G137), .B(KEYINPUT126), .ZN(n764) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(G39) );
endmodule

