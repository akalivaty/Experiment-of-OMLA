//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n546, new_n548, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n459), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT64), .Z(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  INV_X1    g048(.A(new_n462), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n474), .A2(G136), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(G162));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  OAI211_X1 g057(.A(G138), .B(new_n459), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(KEYINPUT4), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT66), .A2(KEYINPUT4), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n461), .A2(G138), .A3(new_n459), .A4(new_n484), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n459), .B2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n481), .C2(new_n482), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT65), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n461), .A2(new_n495), .A3(G126), .A4(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n489), .A2(new_n497), .A3(KEYINPUT67), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n489), .B2(new_n497), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(KEYINPUT68), .A3(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n503), .A2(new_n505), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n512), .B1(G651), .B2(new_n519), .ZN(G166));
  AND2_X1   g095(.A1(new_n506), .A2(new_n507), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n507), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT69), .B(G51), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n508), .A2(new_n534), .B1(new_n510), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n532), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n508), .A2(new_n541), .B1(new_n510), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT70), .Z(G188));
  NOR2_X1   g126(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n510), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OAI221_X1 g131(.A(new_n554), .B1(new_n555), .B2(new_n508), .C1(new_n556), .C2(new_n532), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n558));
  NOR4_X1   g133(.A1(new_n510), .A2(new_n553), .A3(new_n552), .A4(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT72), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(new_n557), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n521), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n523), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND3_X1  g144(.A1(new_n506), .A2(KEYINPUT73), .A3(G61), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n516), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(G86), .B2(new_n521), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n521), .A2(G85), .B1(G47), .B2(new_n523), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n532), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n506), .A2(G92), .A3(new_n507), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G54), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n532), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n584), .B1(new_n591), .B2(G868), .ZN(G284));
  OAI21_X1  g167(.A(new_n584), .B1(new_n591), .B2(G868), .ZN(G321));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G286), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n594), .ZN(G297));
  AOI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n594), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G860), .ZN(G148));
  NOR2_X1   g175(.A1(new_n544), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n591), .A2(new_n599), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT76), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT77), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT11), .Z(G282));
  XOR2_X1   g181(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(G2100), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n608), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n472), .A2(G123), .ZN(new_n612));
  OR2_X1    g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(G111), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n476), .B1(new_n614), .B2(G2105), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n474), .A2(G135), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n612), .A2(G2096), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(G2096), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT79), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT80), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT15), .B(G2435), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT14), .ZN(new_n626));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  AND2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n634), .B2(KEYINPUT81), .ZN(new_n635));
  AOI211_X1 g210(.A(new_n633), .B(new_n635), .C1(KEYINPUT81), .C2(new_n634), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2067), .B(G2678), .Z(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT17), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n640), .B2(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2096), .B(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(G227));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT82), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT19), .Z(new_n652));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n652), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT83), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G23), .ZN(new_n670));
  INV_X1    g245(.A(G288), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT33), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1976), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(G22), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G166), .B2(new_n669), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1971), .ZN(new_n678));
  MUX2_X1   g253(.A(G6), .B(G305), .S(G16), .Z(new_n679));
  XOR2_X1   g254(.A(KEYINPUT32), .B(G1981), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n674), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(KEYINPUT84), .A2(G29), .ZN(new_n686));
  NOR2_X1   g261(.A1(KEYINPUT84), .A2(G29), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G25), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n472), .A2(G119), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  INV_X1    g267(.A(G107), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n476), .B1(new_n693), .B2(G2105), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n474), .A2(G131), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n690), .B1(new_n697), .B2(new_n689), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT35), .B(G1991), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G24), .B(G290), .S(G16), .Z(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(G1986), .Z(new_n703));
  NAND3_X1  g278(.A1(new_n685), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  OR3_X1    g279(.A1(new_n704), .A2(KEYINPUT89), .A3(KEYINPUT36), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT36), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT88), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(KEYINPUT88), .A3(KEYINPUT36), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT89), .B1(new_n704), .B2(KEYINPUT36), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n705), .A2(new_n708), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n591), .A2(new_n669), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G4), .B2(new_n669), .ZN(new_n713));
  INV_X1    g288(.A(G1348), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n669), .A2(G19), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n544), .B2(new_n669), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1341), .Z(new_n719));
  INV_X1    g294(.A(G2084), .ZN(new_n720));
  NAND2_X1  g295(.A1(G160), .A2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G34), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n721), .B1(new_n688), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n472), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT26), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n474), .A2(G141), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n726), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n725), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT27), .B(G1996), .Z(new_n737));
  OAI221_X1 g312(.A(new_n719), .B1(new_n720), .B2(new_n724), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n474), .A2(G139), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT25), .Z(new_n741));
  AOI22_X1  g316(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n741), .C1(new_n459), .C2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT92), .ZN(new_n744));
  MUX2_X1   g319(.A(G33), .B(new_n744), .S(G29), .Z(new_n745));
  AOI211_X1 g320(.A(new_n716), .B(new_n738), .C1(G2072), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G162), .A2(new_n689), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G35), .B2(new_n689), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT98), .B(G1956), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n669), .A2(KEYINPUT23), .A3(G20), .ZN(new_n752));
  AOI21_X1  g327(.A(KEYINPUT23), .B1(new_n669), .B2(G20), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n752), .B(new_n753), .C1(G299), .C2(G16), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n750), .A2(G2090), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n751), .ZN(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n736), .A2(new_n737), .B1(new_n720), .B2(new_n724), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G171), .B2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(G1961), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT97), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n746), .A2(new_n755), .A3(new_n758), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n745), .A2(G2072), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT93), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n669), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n669), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G28), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n771), .B2(KEYINPUT30), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT30), .B2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n612), .A2(new_n616), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n689), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n761), .B2(G1961), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n770), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  AOI21_X1  g354(.A(KEYINPUT28), .B1(new_n689), .B2(G26), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n689), .A2(KEYINPUT28), .A3(G26), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n472), .A2(G128), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n474), .A2(G140), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n459), .A2(G116), .ZN(new_n785));
  OR3_X1    g360(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n786));
  OAI21_X1  g361(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n786), .A2(G2104), .A3(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n788), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n780), .B(new_n782), .C1(new_n789), .C2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT91), .B(G2067), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n766), .A2(new_n779), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n688), .A2(G27), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n688), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2078), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n764), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n711), .A2(new_n715), .A3(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  AOI22_X1  g374(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n532), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  INV_X1    g377(.A(G55), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n508), .A2(new_n802), .B1(new_n510), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT100), .B1(new_n801), .B2(new_n804), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT101), .B(G860), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  AOI21_X1  g387(.A(new_n544), .B1(new_n807), .B2(new_n808), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n805), .A2(new_n540), .A3(new_n543), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT99), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(KEYINPUT99), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n591), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(new_n810), .ZN(G145));
  XNOR2_X1  g397(.A(new_n774), .B(G160), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G162), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n487), .A2(new_n488), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT102), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n825), .B1(new_n830), .B2(new_n497), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT102), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT102), .B1(new_n487), .B2(new_n488), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n825), .B(new_n497), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n789), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n789), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n734), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n735), .A3(new_n838), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n840), .A2(new_n743), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n744), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n472), .A2(G130), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n474), .A2(G142), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n459), .A2(G118), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n476), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI221_X1 g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .C1(G106), .C2(G2105), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n844), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n610), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n696), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n842), .A2(new_n843), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n840), .A2(new_n841), .ZN(new_n855));
  INV_X1    g430(.A(new_n744), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n840), .A2(new_n743), .A3(new_n841), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n824), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n852), .B1(new_n842), .B2(new_n843), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(new_n854), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(KEYINPUT105), .A3(new_n824), .ZN(new_n866));
  AOI21_X1  g441(.A(G37), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  INV_X1    g443(.A(new_n824), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT105), .B1(new_n865), .B2(new_n824), .ZN(new_n873));
  AOI211_X1 g448(.A(new_n861), .B(new_n869), .C1(new_n863), .C2(new_n864), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n872), .B(new_n870), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT106), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT40), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT40), .B1(new_n871), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(G395));
  NAND2_X1  g454(.A1(new_n809), .A2(new_n594), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n817), .B(new_n602), .Z(new_n881));
  NAND2_X1  g456(.A1(G299), .A2(new_n590), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n591), .A2(new_n561), .A3(new_n563), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n882), .B2(new_n883), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(new_n881), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(G305), .B(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G166), .ZN(new_n892));
  XOR2_X1   g467(.A(G290), .B(KEYINPUT107), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n890), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n880), .B1(new_n896), .B2(new_n594), .ZN(G295));
  OAI21_X1  g472(.A(new_n880), .B1(new_n896), .B2(new_n594), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n899));
  XNOR2_X1  g474(.A(G301), .B(G286), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n817), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n815), .A2(new_n816), .A3(new_n900), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n815), .A2(KEYINPUT108), .A3(new_n816), .A4(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n888), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n884), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n902), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n899), .B1(new_n895), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n894), .A2(KEYINPUT109), .A3(new_n907), .A4(new_n909), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n872), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n884), .B1(new_n905), .B2(new_n906), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT110), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n902), .A2(new_n904), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n888), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n894), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n911), .B2(new_n912), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n916), .A2(new_n918), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n894), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n895), .A2(new_n910), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n922), .A2(new_n926), .A3(new_n929), .A4(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n925), .B2(KEYINPUT43), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n934), .ZN(G397));
  XOR2_X1   g510(.A(new_n789), .B(G2067), .Z(new_n936));
  NAND2_X1  g511(.A1(new_n734), .A2(G1996), .ZN(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n735), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n697), .A2(new_n700), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n696), .A2(new_n699), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT112), .B1(new_n836), .B2(G1384), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n497), .B1(new_n832), .B2(new_n833), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT103), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n834), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G160), .A2(G40), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n946), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g535(.A1(G286), .A2(G8), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT119), .Z(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT67), .ZN(new_n964));
  INV_X1    g539(.A(new_n492), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n495), .B1(new_n471), .B2(G126), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n493), .A2(KEYINPUT65), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n968), .B2(new_n826), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n489), .A2(new_n497), .A3(KEYINPUT67), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n953), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(new_n956), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n830), .B2(new_n497), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AND4_X1   g551(.A1(new_n720), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n949), .A2(new_n953), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n956), .B1(new_n978), .B2(new_n948), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n953), .A4(new_n970), .ZN(new_n980));
  AOI21_X1  g555(.A(G1966), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n963), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n973), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n984));
  INV_X1    g559(.A(new_n980), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n769), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n972), .A2(new_n976), .A3(new_n720), .A4(new_n973), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n982), .B(KEYINPUT51), .C1(new_n963), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT120), .ZN(new_n990));
  OAI21_X1  g565(.A(G8), .B1(new_n977), .B2(new_n981), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n962), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n990), .B1(new_n989), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n960), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n982), .A2(KEYINPUT51), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n988), .A2(new_n963), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT120), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(KEYINPUT62), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n953), .C1(new_n831), .C2(new_n835), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n956), .B1(new_n971), .B2(new_n948), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(G2078), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n956), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n976), .ZN(new_n1009));
  INV_X1    g584(.A(G1961), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G2078), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n979), .A2(new_n1013), .A3(new_n980), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n979), .A2(KEYINPUT121), .A3(new_n1013), .A4(new_n980), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n978), .A2(new_n956), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n983), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1023), .C1(new_n1022), .C2(G288), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G305), .A2(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n576), .A2(new_n1026), .A3(new_n578), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1021), .A3(new_n1031), .ZN(new_n1032));
  OAI221_X1 g607(.A(G8), .B1(new_n1022), .B2(G288), .C1(new_n978), .C2(new_n956), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1033), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n1033), .B2(KEYINPUT52), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1024), .B(new_n1032), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G166), .A2(new_n983), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1008), .A2(new_n757), .A3(new_n976), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1971), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1042));
  OAI211_X1 g617(.A(G8), .B(new_n1039), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n500), .A2(KEYINPUT114), .A3(new_n975), .A4(new_n953), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n969), .A2(new_n975), .A3(new_n953), .A4(new_n970), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n956), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n757), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1006), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n983), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1037), .B(new_n1043), .C1(new_n1039), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n996), .A2(new_n1002), .A3(new_n1019), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1032), .A2(new_n1022), .A3(new_n671), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1027), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1021), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1043), .B2(new_n1036), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n983), .B1(new_n1052), .B2(new_n1040), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1037), .B(new_n1061), .C1(new_n1039), .C2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1039), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n1064), .B2(new_n1036), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n988), .A2(G168), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1039), .B2(new_n1062), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1063), .A2(new_n1065), .A3(KEYINPUT63), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT63), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1054), .B2(new_n1066), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1060), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1056), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(new_n973), .A3(new_n1049), .ZN(new_n1074));
  INV_X1    g649(.A(G1956), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n560), .B(KEYINPUT57), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1004), .A2(new_n1005), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1004), .A2(new_n1005), .A3(new_n1082), .A4(new_n1079), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1076), .A2(new_n1078), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1020), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(G2067), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1348), .B1(new_n1008), .B2(new_n976), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1084), .B(new_n591), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1956), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1077), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1084), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1006), .A2(G1996), .B1(new_n1020), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n544), .A2(KEYINPUT117), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1091), .A2(new_n1084), .A3(KEYINPUT61), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1096), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1087), .A2(new_n1086), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT118), .A3(new_n591), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT118), .B1(new_n1111), .B2(new_n591), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1093), .B1(new_n1107), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n952), .B1(new_n951), .B2(new_n953), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT112), .B(G1384), .C1(new_n950), .C2(new_n834), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1120), .A2(new_n1121), .A3(KEYINPUT45), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT122), .B1(new_n1122), .B2(new_n956), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1004), .A2(new_n1013), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n955), .A2(new_n1125), .A3(new_n973), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(KEYINPUT53), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(G301), .A3(new_n1012), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1019), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n994), .A2(new_n1054), .A3(new_n995), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1012), .A2(new_n1134), .A3(G301), .A4(new_n1018), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1018), .A2(G301), .A3(new_n1007), .A4(new_n1011), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1131), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1127), .A2(new_n1012), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(G301), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1119), .A2(new_n1132), .A3(new_n1133), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n959), .B1(new_n1072), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n957), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n944), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT48), .Z(new_n1145));
  NOR2_X1   g720(.A1(new_n943), .A2(new_n1143), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT126), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1143), .B2(G1996), .ZN(new_n1150));
  INV_X1    g725(.A(new_n936), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n957), .B1(new_n734), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n957), .B(new_n938), .C1(new_n1153), .C2(KEYINPUT46), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT47), .ZN(new_n1156));
  INV_X1    g731(.A(new_n942), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n940), .A2(new_n1157), .B1(G2067), .B2(new_n789), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n957), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT124), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1148), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n1142), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1132), .A2(new_n1140), .A3(new_n1133), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1091), .A2(new_n1084), .A3(KEYINPUT61), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT61), .B1(new_n1091), .B2(new_n1084), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1104), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1092), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1056), .A2(new_n1071), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n958), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1161), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1162), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g750(.A1(new_n871), .A2(new_n876), .ZN(new_n1177));
  INV_X1    g751(.A(G319), .ZN(new_n1178));
  NOR2_X1   g752(.A1(G229), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g753(.A1(G401), .A2(G227), .ZN(new_n1180));
  AND4_X1   g754(.A1(new_n1177), .A2(new_n932), .A3(new_n1179), .A4(new_n1180), .ZN(G308));
  NAND4_X1  g755(.A1(new_n1177), .A2(new_n932), .A3(new_n1179), .A4(new_n1180), .ZN(G225));
endmodule


