//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(G222), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n247), .B(new_n248), .C1(new_n249), .C2(new_n245), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(new_n252), .A3(G274), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n252), .A2(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(G226), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G179), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n216), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n206), .A2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n268), .A2(new_n270), .B1(G50), .B2(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(G58), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT8), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT67), .B1(new_n277), .B2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(new_n207), .A3(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n266), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(G169), .B1(new_n254), .B2(new_n261), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n263), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G244), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n257), .B1(new_n288), .B2(new_n259), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n245), .A2(G232), .A3(new_n246), .ZN(new_n291));
  INV_X1    g0091(.A(G107), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n290), .B(new_n291), .C1(new_n292), .C2(new_n245), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n289), .B1(new_n293), .B2(new_n253), .ZN(new_n294));
  INV_X1    g0094(.A(G200), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n207), .A2(new_n277), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT68), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT68), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n276), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G20), .A2(G77), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(KEYINPUT69), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n207), .A2(G33), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT69), .B1(new_n301), .B2(new_n302), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n265), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n267), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  INV_X1    g0111(.A(new_n267), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n265), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n313), .A3(G77), .A4(new_n269), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n249), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n294), .A2(G190), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n296), .A2(new_n309), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n309), .A2(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n294), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G169), .B2(new_n294), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n318), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n295), .B1(new_n254), .B2(new_n261), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n285), .B2(KEYINPUT9), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT9), .ZN(new_n330));
  NOR4_X1   g0130(.A1(new_n271), .A2(new_n284), .A3(KEYINPUT71), .A4(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n327), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n254), .A2(new_n261), .A3(G190), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n330), .B1(new_n271), .B2(new_n284), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(new_n325), .C2(new_n326), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT10), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n326), .B1(new_n262), .B2(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n334), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n285), .A2(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT71), .ZN(new_n341));
  INV_X1    g0141(.A(new_n331), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT10), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .A4(new_n327), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n287), .B(new_n324), .C1(new_n336), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G68), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n272), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n348), .B2(new_n201), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n282), .A2(G159), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NOR4_X1   g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .A4(G20), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n353), .B2(new_n354), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n277), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(KEYINPUT77), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n362), .A3(new_n207), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n356), .B1(new_n363), .B2(new_n355), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT16), .B(new_n352), .C1(new_n364), .C2(new_n347), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n355), .B1(new_n245), .B2(G20), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n353), .A2(new_n354), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n347), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n366), .B1(new_n370), .B2(new_n351), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n365), .A2(new_n265), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n276), .A2(new_n269), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n268), .A2(new_n373), .B1(new_n267), .B2(new_n276), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT78), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n368), .B2(new_n207), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n378), .B2(new_n356), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n352), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n266), .B1(new_n380), .B2(new_n366), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n374), .B1(new_n381), .B2(new_n365), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT78), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT18), .ZN(new_n385));
  OAI211_X1 g0185(.A(G226), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT79), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT79), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n245), .A2(new_n388), .A3(G226), .A4(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(G223), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n252), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G232), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n257), .B1(new_n396), .B2(new_n259), .ZN(new_n397));
  OAI21_X1  g0197(.A(G169), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n397), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n393), .B1(new_n389), .B2(new_n387), .ZN(new_n400));
  OAI211_X1 g0200(.A(G179), .B(new_n399), .C1(new_n400), .C2(new_n252), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n377), .A2(new_n384), .A3(new_n385), .A4(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(G190), .B(new_n399), .C1(new_n400), .C2(new_n252), .ZN(new_n404));
  OAI21_X1  g0204(.A(G200), .B1(new_n395), .B2(new_n397), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n372), .A2(new_n375), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n382), .A2(KEYINPUT17), .A3(new_n404), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n377), .A2(new_n384), .A3(new_n402), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(KEYINPUT18), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n346), .A2(new_n403), .A3(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(G226), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n245), .A2(KEYINPUT73), .A3(G226), .A4(new_n246), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n245), .A2(G232), .A3(G1698), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n253), .ZN(new_n421));
  INV_X1    g0221(.A(G238), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n257), .B1(new_n422), .B2(new_n259), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT74), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n420), .B2(new_n253), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n427), .A3(KEYINPUT13), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(G169), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n431), .A2(new_n435), .A3(G169), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n428), .A2(new_n429), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n426), .A2(G179), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n278), .A2(new_n280), .A3(G77), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n207), .B2(G68), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n441), .A2(KEYINPUT75), .B1(new_n202), .B2(new_n297), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n265), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT11), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n312), .A2(new_n347), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT12), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n310), .A2(new_n313), .A3(G68), .A4(new_n269), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT76), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n449), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(KEYINPUT11), .B(new_n265), .C1(new_n442), .C2(new_n443), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n446), .A2(new_n450), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n439), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n426), .A2(G190), .A3(new_n437), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n455), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n431), .A2(G200), .A3(new_n432), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n413), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT89), .ZN(new_n463));
  OAI211_X1 g0263(.A(G257), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n464));
  OAI211_X1 g0264(.A(G250), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G294), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  INV_X1    g0270(.A(new_n216), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n468), .A2(new_n470), .B1(new_n471), .B2(new_n251), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n467), .A2(new_n253), .B1(new_n472), .B2(G264), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n468), .A2(G274), .A3(new_n252), .A4(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(G179), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G169), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n463), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n478), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(KEYINPUT89), .A3(new_n475), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n207), .B(G87), .C1(new_n353), .C2(new_n354), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n245), .A2(new_n484), .A3(new_n207), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G116), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT23), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n207), .B2(G107), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n292), .A2(KEYINPUT23), .A3(G20), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n486), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n487), .B1(new_n486), .B2(new_n493), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n265), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n312), .A2(new_n292), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n206), .A2(G33), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n266), .A2(new_n499), .A3(new_n267), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n267), .A2(new_n500), .A3(new_n216), .A4(new_n264), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n498), .B1(G107), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n479), .A2(new_n481), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n473), .A2(new_n474), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n473), .A2(G190), .A3(new_n474), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n496), .A2(new_n509), .A3(new_n505), .A4(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G238), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n488), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n253), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT83), .B1(new_n469), .B2(G1), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT83), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n206), .A3(G45), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n252), .A2(new_n517), .A3(new_n519), .A4(G250), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n252), .A2(G274), .A3(new_n470), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT84), .B1(new_n524), .B2(G179), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n253), .B2(new_n515), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT84), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n321), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT85), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT85), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G87), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n207), .B1(new_n418), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n245), .A2(new_n207), .A3(G68), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n536), .B1(new_n305), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n265), .B1(new_n312), .B2(new_n304), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT87), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT86), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n304), .B(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n504), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n504), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n524), .A2(new_n477), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n529), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n504), .A2(G87), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n543), .B(new_n552), .C1(new_n295), .C2(new_n526), .ZN(new_n553));
  INV_X1    g0353(.A(G190), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n524), .A2(new_n554), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G13), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(G1), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(G20), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n264), .A2(new_n216), .B1(G20), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(new_n207), .C1(G33), .C2(new_n540), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT20), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n560), .B1(new_n206), .B2(G33), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n310), .A2(new_n313), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT5), .A2(G41), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT5), .A2(G41), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n470), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(G270), .A3(new_n252), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n474), .ZN(new_n575));
  OAI211_X1 g0375(.A(G264), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n576));
  OAI211_X1 g0376(.A(G257), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n245), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n253), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n570), .B(KEYINPUT88), .C1(new_n580), .C2(new_n295), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT88), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n574), .A2(new_n474), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n253), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n295), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n310), .A2(new_n313), .A3(new_n568), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n561), .C1(new_n566), .C2(new_n565), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n582), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n580), .A2(G190), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n581), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(new_n584), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT21), .A4(G169), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n580), .A3(G179), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n591), .A3(G169), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  AND2_X1   g0399(.A1(G97), .A2(G107), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n534), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT6), .A2(G97), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT80), .B1(new_n602), .B2(G107), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(new_n292), .A3(KEYINPUT6), .A4(G97), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n607));
  OAI21_X1  g0407(.A(G107), .B1(new_n378), .B2(new_n356), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n265), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n267), .A2(G97), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n504), .B2(G97), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n573), .A2(G257), .A3(new_n252), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n474), .ZN(new_n614));
  OAI211_X1 g0414(.A(G244), .B(new_n246), .C1(new_n353), .C2(new_n354), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT4), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n245), .A2(G244), .A3(new_n246), .A4(new_n617), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n245), .A2(G250), .A3(G1698), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .A4(new_n563), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n622), .B2(new_n253), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n610), .B(new_n612), .C1(new_n295), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(G190), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n504), .A2(G97), .ZN(new_n627));
  INV_X1    g0427(.A(new_n611), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n266), .B1(new_n607), .B2(new_n608), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n623), .B2(G169), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n622), .A2(new_n253), .ZN(new_n632));
  INV_X1    g0432(.A(new_n614), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G179), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n624), .A2(new_n626), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n598), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n462), .A2(new_n512), .A3(new_n557), .A4(new_n637), .ZN(G372));
  AOI21_X1  g0438(.A(new_n555), .B1(new_n553), .B2(KEYINPUT90), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n524), .A2(G200), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT90), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n543), .A4(new_n552), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n526), .A2(new_n321), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n550), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n639), .A2(new_n642), .B1(new_n549), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n631), .A2(new_n635), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT26), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(KEYINPUT26), .A2(new_n646), .A3(new_n551), .A4(new_n556), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n549), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n634), .A2(G200), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n610), .A3(new_n612), .A4(new_n625), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n610), .A2(new_n612), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n623), .A2(new_n321), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(new_n654), .C1(G169), .C2(new_n623), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n597), .A2(new_n593), .A3(new_n592), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n496), .A2(new_n505), .B1(new_n480), .B2(new_n475), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n652), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n543), .A2(new_n552), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n526), .A2(new_n295), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT90), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n555), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n642), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n511), .A3(new_n650), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n650), .B1(new_n658), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n462), .B1(new_n649), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n376), .A2(new_n402), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT18), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n376), .A2(new_n385), .A3(new_n402), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n320), .A2(new_n323), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n439), .A2(new_n455), .B1(new_n460), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n672), .B2(new_n410), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n336), .A2(new_n345), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n287), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n666), .A2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n507), .A2(new_n511), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n559), .A2(new_n207), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n559), .A2(new_n680), .A3(new_n207), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT91), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n679), .A2(KEYINPUT91), .A3(G213), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n656), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n506), .B1(new_n478), .B2(new_n476), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n677), .A2(new_n690), .B1(new_n691), .B2(new_n688), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT92), .ZN(new_n693));
  INV_X1    g0493(.A(new_n506), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n512), .B1(new_n694), .B2(new_n689), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n507), .A2(new_n689), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n689), .A2(new_n570), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n656), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n598), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n693), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n210), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n535), .A2(G116), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n708), .A3(new_n206), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(KEYINPUT93), .B1(new_n215), .B2(new_n706), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(KEYINPUT93), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n663), .A2(KEYINPUT26), .A3(new_n646), .A4(new_n650), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT95), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT26), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n551), .A2(new_n556), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n655), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n663), .A2(new_n511), .A3(new_n650), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n597), .A2(new_n593), .A3(new_n592), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n507), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT96), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n636), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n655), .A2(KEYINPUT96), .A3(new_n652), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n721), .A2(new_n723), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n650), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT29), .B(new_n689), .C1(new_n720), .C2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n689), .B1(new_n649), .B2(new_n665), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n688), .A2(KEYINPUT31), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n583), .A2(new_n584), .A3(G179), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n526), .A2(new_n473), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT30), .A4(new_n623), .ZN(new_n739));
  AOI21_X1  g0539(.A(G179), .B1(new_n583), .B2(new_n584), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n634), .A2(new_n740), .A3(new_n508), .A4(new_n524), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n632), .A2(new_n526), .A3(new_n473), .A4(new_n633), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(new_n736), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n735), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT94), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n748), .B(new_n743), .C1(new_n744), .C2(new_n736), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n747), .A2(new_n749), .A3(new_n739), .A4(new_n741), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n688), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n637), .A2(new_n512), .A3(new_n557), .A4(new_n689), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n734), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n733), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n712), .B1(new_n758), .B2(G1), .ZN(G364));
  INV_X1    g0559(.A(new_n706), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n558), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n206), .B1(new_n761), .B2(G45), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n700), .A2(G330), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n702), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n700), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n763), .B(KEYINPUT97), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n216), .B1(G20), .B2(new_n477), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n776), .A2(new_n207), .A3(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT32), .Z(new_n779));
  OAI21_X1  g0579(.A(G20), .B1(new_n776), .B2(new_n554), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G97), .ZN(new_n781));
  NAND2_X1  g0581(.A1(G20), .A2(G179), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n782), .A2(new_n295), .A3(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n245), .B1(new_n784), .B2(new_n249), .C1(new_n347), .C2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n531), .A2(new_n533), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n207), .A2(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(new_n554), .A3(G200), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n788), .A2(new_n790), .B1(new_n791), .B2(new_n292), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n782), .A2(new_n554), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n782), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(G190), .A3(G200), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n794), .A2(new_n272), .B1(new_n796), .B2(new_n202), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n787), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n779), .A2(new_n781), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G326), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n802), .A2(new_n791), .B1(new_n790), .B2(new_n578), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G322), .C2(new_n793), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n780), .A2(G294), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n777), .A2(G329), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n784), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n245), .B(new_n808), .C1(new_n785), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n774), .B1(new_n799), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n243), .A2(new_n469), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n358), .A2(new_n362), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n705), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n469), .B2(new_n215), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n813), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n705), .A2(new_n368), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n822), .A2(G355), .B1(new_n560), .B2(new_n705), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n768), .A2(new_n773), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n772), .B(new_n812), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n765), .B1(new_n770), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  OAI221_X1 g0628(.A(new_n368), .B1(new_n790), .B2(new_n292), .C1(new_n784), .C2(new_n560), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n786), .A2(KEYINPUT100), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n829), .B1(new_n833), .B2(G283), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n777), .A2(G311), .ZN(new_n835));
  INV_X1    g0635(.A(G294), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n794), .A2(new_n836), .B1(new_n796), .B2(new_n578), .ZN(new_n837));
  INV_X1    g0637(.A(new_n791), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(G87), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n834), .A2(new_n781), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G150), .A2(new_n785), .B1(new_n783), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n796), .C1(new_n843), .C2(new_n794), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT34), .Z(new_n845));
  NOR2_X1   g0645(.A1(new_n791), .A2(new_n347), .ZN(new_n846));
  INV_X1    g0646(.A(new_n790), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n846), .B(new_n814), .C1(G50), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n780), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  INV_X1    g0650(.A(new_n777), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n848), .B1(new_n272), .B2(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n840), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n854), .A2(new_n855), .A3(new_n774), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n773), .A2(new_n766), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n772), .B(new_n856), .C1(new_n249), .C2(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT102), .Z(new_n859));
  NAND2_X1  g0659(.A1(new_n319), .A2(new_n688), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT103), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n319), .A2(new_n862), .A3(new_n688), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n318), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n320), .A2(new_n323), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n671), .A2(new_n689), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n859), .B1(new_n766), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n730), .A2(new_n868), .ZN(new_n870));
  INV_X1    g0670(.A(new_n867), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n864), .B2(new_n865), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n872), .B(new_n689), .C1(new_n649), .C2(new_n665), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n870), .A2(new_n755), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n763), .B1(new_n875), .B2(new_n756), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n869), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(G384));
  NOR2_X1   g0678(.A1(new_n761), .A2(new_n206), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n411), .A2(KEYINPUT18), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n408), .A2(new_n409), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n403), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n365), .A2(new_n265), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n352), .B1(new_n364), .B2(new_n347), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n366), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n374), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n686), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n406), .B1(new_n887), .B2(new_n686), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n398), .A2(new_n401), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n686), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n377), .A2(new_n384), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n406), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n411), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n893), .B2(new_n898), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n900), .A2(new_n901), .B1(new_n889), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT31), .B1(new_n750), .B2(new_n688), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n868), .B1(new_n906), .B2(new_n754), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n455), .A2(new_n688), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n456), .A2(new_n460), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n460), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n455), .B(new_n688), .C1(new_n910), .C2(new_n439), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n880), .B1(new_n903), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n899), .A2(KEYINPUT38), .ZN(new_n915));
  INV_X1    g0715(.A(new_n888), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n412), .B2(new_n403), .ZN(new_n917));
  AOI211_X1 g0717(.A(KEYINPUT78), .B(new_n374), .C1(new_n381), .C2(new_n365), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n383), .B1(new_n372), .B2(new_n375), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n918), .A2(new_n919), .A3(new_n686), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n667), .A2(new_n406), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n668), .A2(new_n408), .A3(new_n409), .A4(new_n669), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n898), .B1(new_n923), .B2(new_n920), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n915), .A2(new_n917), .B1(new_n924), .B2(KEYINPUT38), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n925), .A2(KEYINPUT40), .A3(new_n912), .A4(new_n907), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n751), .A2(new_n752), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n754), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n462), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n734), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n925), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n439), .A2(new_n455), .A3(new_n689), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n889), .A2(new_n902), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n883), .A2(new_n888), .B1(new_n893), .B2(new_n898), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n938), .B(KEYINPUT39), .C1(KEYINPUT38), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n670), .A2(new_n894), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n873), .A2(new_n867), .B1(new_n909), .B2(new_n911), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n938), .B1(new_n939), .B2(KEYINPUT38), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n729), .A2(new_n462), .A3(new_n732), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n675), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n879), .B1(new_n933), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n933), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(G116), .A3(new_n217), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n214), .A2(new_n249), .A3(new_n348), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n347), .A2(G50), .ZN(new_n957));
  OAI211_X1 g0757(.A(G1), .B(new_n558), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(G367));
  NOR2_X1   g0759(.A1(new_n655), .A2(new_n689), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT104), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n653), .A2(new_n688), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n725), .A2(new_n726), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n655), .B1(new_n965), .B2(new_n507), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n689), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n677), .A2(new_n690), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT42), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n965), .A2(KEYINPUT42), .A3(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n688), .A2(new_n659), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n645), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n650), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT105), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n703), .A2(new_n965), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n976), .B1(new_n971), .B2(new_n978), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n706), .B(KEYINPUT41), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n693), .A2(new_n964), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n693), .A2(new_n990), .A3(new_n964), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n693), .B2(new_n964), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n703), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n695), .A2(new_n696), .A3(new_n690), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT106), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n695), .A2(KEYINPUT106), .A3(new_n696), .A4(new_n690), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n968), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(new_n702), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n989), .A2(new_n993), .A3(new_n703), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n996), .A2(new_n758), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n986), .B1(new_n1004), .B2(new_n758), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n762), .B(KEYINPUT107), .Z(new_n1006));
  OAI211_X1 g0806(.A(new_n984), .B(new_n985), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT109), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n825), .B1(new_n210), .B2(new_n304), .C1(new_n817), .C2(new_n235), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n245), .B1(new_n790), .B2(new_n272), .C1(new_n784), .C2(new_n202), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n833), .B2(G159), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n780), .A2(G68), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n796), .A2(new_n843), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n791), .A2(new_n249), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G150), .C2(new_n793), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n777), .A2(G137), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n815), .B1(G283), .B2(new_n783), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n836), .B2(new_n832), .C1(new_n1019), .C2(new_n851), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n847), .A2(G116), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT46), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n796), .A2(new_n807), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n791), .A2(new_n540), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G303), .C2(new_n793), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1022), .B(new_n1025), .C1(new_n292), .C2(new_n849), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1017), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT47), .Z(new_n1028));
  OAI211_X1 g0828(.A(new_n771), .B(new_n1009), .C1(new_n1028), .C2(new_n774), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT108), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n769), .B2(new_n974), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1007), .A2(new_n1008), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1008), .B1(new_n1007), .B2(new_n1031), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(G387));
  NOR2_X1   g0835(.A1(new_n697), .A2(new_n769), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n708), .C1(G68), .C2(G77), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n276), .A2(new_n202), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n817), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT110), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1041), .A2(new_n1042), .B1(G45), .B2(new_n232), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n822), .A2(new_n708), .B1(new_n292), .B2(new_n705), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n825), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n771), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n794), .A2(new_n202), .B1(new_n790), .B2(new_n249), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n796), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1024), .B(new_n1049), .C1(G159), .C2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n784), .A2(new_n347), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n814), .B(new_n1052), .C1(new_n276), .C2(new_n785), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n780), .A2(new_n546), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT111), .B(G150), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n777), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n833), .A2(G311), .B1(G322), .B2(new_n1050), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G303), .A2(new_n783), .B1(new_n793), .B2(G317), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT48), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n849), .A2(new_n802), .B1(new_n836), .B2(new_n790), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n815), .B1(G116), .B2(new_n838), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n800), .C2(new_n851), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT49), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1057), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1036), .B(new_n1048), .C1(new_n1071), .C2(new_n773), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1002), .A2(new_n758), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n706), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1002), .A2(new_n758), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(new_n1003), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n703), .B1(new_n989), .B2(new_n993), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1080), .A2(new_n1004), .A3(new_n706), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1006), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n240), .A2(new_n817), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n825), .B1(new_n540), .B2(new_n210), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n771), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n833), .A2(G50), .B1(G143), .B2(new_n777), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n347), .A2(new_n790), .B1(new_n791), .B2(new_n530), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n814), .B(new_n1088), .C1(new_n276), .C2(new_n783), .ZN(new_n1089));
  INV_X1    g0889(.A(G159), .ZN(new_n1090));
  INV_X1    g0890(.A(G150), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n794), .A2(new_n1090), .B1(new_n796), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n780), .A2(G77), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1087), .A2(new_n1089), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n777), .A2(G322), .B1(G283), .B2(new_n847), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT114), .Z(new_n1097));
  OAI221_X1 g0897(.A(new_n368), .B1(new_n791), .B2(new_n292), .C1(new_n784), .C2(new_n836), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n833), .B2(G303), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n794), .A2(new_n807), .B1(new_n796), .B2(new_n1019), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1099), .B(new_n1102), .C1(new_n560), .C2(new_n849), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1095), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1086), .B1(new_n1104), .B2(new_n773), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n964), .B2(new_n769), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1081), .A2(new_n1083), .A3(new_n1106), .ZN(G390));
  AND2_X1   g0907(.A1(new_n909), .A2(new_n911), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n930), .A2(G330), .A3(new_n872), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n873), .A2(new_n867), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n912), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n935), .A2(new_n940), .B1(new_n1112), .B2(new_n936), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n689), .B(new_n866), .C1(new_n720), .C2(new_n728), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1114), .A2(new_n867), .B1(new_n909), .B2(new_n911), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n925), .A2(new_n936), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1110), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n636), .B1(new_n722), .B2(new_n691), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1119), .A2(new_n721), .B1(new_n549), .B2(new_n644), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n557), .A2(KEYINPUT26), .A3(new_n646), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n663), .A2(new_n650), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n716), .B1(new_n1122), .B2(new_n655), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n688), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n871), .B1(new_n1125), .B2(new_n872), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n936), .B1(new_n1126), .B2(new_n1108), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n940), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n923), .A2(new_n920), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n411), .A2(new_n895), .A3(new_n897), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n667), .A2(new_n406), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n896), .B1(new_n1131), .B2(new_n895), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n901), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT39), .B1(new_n1134), .B2(new_n938), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1127), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1114), .A2(new_n867), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n912), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n937), .B1(new_n1134), .B2(new_n938), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n734), .B(new_n868), .C1(new_n753), .C2(new_n754), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n912), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1118), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n912), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1111), .B1(new_n1110), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n1142), .A3(new_n867), .A4(new_n1114), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n462), .A2(G330), .A3(new_n930), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n947), .A2(new_n1150), .A3(new_n675), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1144), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1118), .A2(new_n1143), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n706), .A3(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1118), .A2(new_n1143), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n766), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n857), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n771), .B1(new_n276), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT115), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n245), .B(new_n846), .C1(G97), .C2(new_n783), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n292), .B2(new_n832), .C1(new_n836), .C2(new_n851), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G87), .A2(new_n847), .B1(new_n1050), .B2(G283), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1094), .B(new_n1165), .C1(new_n560), .C2(new_n794), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n847), .A2(new_n1055), .ZN(new_n1167));
  XOR2_X1   g0967(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1168));
  AOI22_X1  g0968(.A1(new_n777), .A2(G125), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n842), .B2(new_n832), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n780), .A2(G159), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n838), .A2(G50), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT54), .B(G143), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n368), .B1(new_n1174), .B2(new_n783), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1050), .A2(G128), .B1(G132), .B2(new_n793), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1164), .A2(new_n1166), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1162), .B1(new_n773), .B2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1158), .A2(new_n1006), .B1(new_n1159), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1157), .A2(new_n1180), .ZN(G378));
  AND2_X1   g0981(.A1(new_n907), .A2(new_n912), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n880), .B1(new_n1134), .B2(new_n938), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n734), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n287), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n285), .B(new_n686), .C1(new_n674), .C2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n686), .A2(new_n285), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n287), .B(new_n1187), .C1(new_n336), .C2(new_n345), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OR3_X1    g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1184), .A2(new_n914), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1184), .B2(new_n914), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n946), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n941), .A2(new_n945), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1193), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n926), .A2(G330), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT40), .B1(new_n1182), .B2(new_n944), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1184), .A2(new_n914), .A3(new_n1193), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1006), .B1(new_n1196), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1198), .A2(new_n766), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n763), .B1(G50), .B2(new_n1160), .ZN(new_n1206));
  INV_X1    g1006(.A(G41), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n814), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT117), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n272), .A2(new_n791), .B1(new_n790), .B2(new_n249), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1211), .B(new_n1208), .C1(G283), .C2(new_n777), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT118), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n546), .A2(new_n783), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n786), .A2(new_n540), .B1(new_n796), .B2(new_n560), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G107), .B2(new_n793), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1012), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1210), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n794), .A2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n786), .A2(new_n850), .B1(new_n784), .B2(new_n842), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G125), .C2(new_n1050), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n847), .A2(new_n1174), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT119), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(new_n1091), .C2(new_n849), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n838), .C2(G159), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(KEYINPUT120), .B(G124), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1229), .C1(new_n851), .C2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1219), .B1(new_n1218), .B2(new_n1217), .C1(new_n1227), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1206), .B1(new_n1232), .B2(new_n773), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1205), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1204), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n946), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1201), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n760), .B1(new_n1243), .B2(new_n1239), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1235), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n1108), .A2(new_n766), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n771), .B1(G68), .B2(new_n1160), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n245), .B(new_n1014), .C1(G107), .C2(new_n783), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n560), .B2(new_n832), .C1(new_n578), .C2(new_n851), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G97), .A2(new_n847), .B1(new_n1050), .B2(G294), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1054), .B(new_n1251), .C1(new_n802), .C2(new_n794), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n814), .B1(G150), .B2(new_n783), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n832), .B2(new_n1173), .C1(new_n1220), .C2(new_n851), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n847), .A2(G159), .B1(new_n838), .B2(G58), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1050), .A2(G132), .B1(G137), .B2(new_n793), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n849), .C2(new_n202), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1250), .A2(new_n1252), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1248), .B1(new_n1258), .B2(new_n773), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1149), .A2(new_n1006), .B1(new_n1247), .B2(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1155), .A2(new_n986), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(G381));
  OR2_X1    g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(G390), .A2(new_n1264), .A3(G384), .A4(G381), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1034), .A2(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1266), .A2(KEYINPUT121), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(KEYINPUT121), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(G375), .A2(G378), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(G407));
  INV_X1    g1070(.A(G213), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1269), .B2(new_n687), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G407), .A2(new_n1272), .ZN(G409));
  NOR3_X1   g1073(.A1(new_n1032), .A2(new_n1033), .A3(G390), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1007), .A2(new_n1031), .A3(G390), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1264), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1007), .A2(new_n1279), .A3(new_n1031), .A4(G390), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1276), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1275), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G390), .B1(new_n1007), .B2(new_n1031), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1278), .A2(KEYINPUT124), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1278), .A2(KEYINPUT124), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1274), .A2(new_n1281), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1271), .A2(G343), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1238), .A2(new_n1006), .B1(new_n1205), .B2(new_n1233), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1203), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n706), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G378), .B(new_n1292), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT122), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1300), .A2(KEYINPUT122), .A3(G378), .A4(new_n1292), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1240), .A2(new_n986), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G378), .B1(new_n1303), .B2(new_n1292), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1291), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1262), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n706), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1260), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n877), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1310), .A2(G384), .A3(new_n1260), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1291), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1314), .B(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1304), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1318), .A2(new_n1291), .A3(new_n1314), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  OAI221_X1 g1120(.A(new_n1290), .B1(new_n1306), .B2(new_n1317), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1289), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1301), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT122), .B1(new_n1245), .B2(G378), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1305), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1327), .A2(KEYINPUT63), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1291), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1326), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1288), .ZN(new_n1331));
  XOR2_X1   g1131(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1306), .B2(new_n1327), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1290), .B1(new_n1306), .B2(new_n1317), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT126), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1330), .B(new_n1288), .C1(new_n1319), .C2(new_n1332), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT126), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1338), .A2(new_n1339), .A3(new_n1335), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1323), .B1(new_n1337), .B2(new_n1340), .ZN(G405));
  OAI22_X1  g1141(.A1(new_n1324), .A2(new_n1325), .B1(G378), .B2(new_n1245), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT127), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1342), .A2(KEYINPUT127), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1327), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  OR2_X1    g1146(.A1(new_n1342), .A2(KEYINPUT127), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1314), .A3(new_n1343), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1346), .A2(new_n1348), .A3(new_n1289), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1289), .B1(new_n1346), .B2(new_n1348), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(G402));
endmodule


