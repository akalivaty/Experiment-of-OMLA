

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G1966), .A2(n826), .ZN(n747) );
  NOR2_X1 U554 ( .A1(KEYINPUT33), .A2(n762), .ZN(n764) );
  NOR2_X2 U555 ( .A1(n759), .A2(n826), .ZN(n760) );
  NAND2_X2 U556 ( .A1(n732), .A2(G8), .ZN(n826) );
  NOR2_X1 U557 ( .A1(n692), .A2(n691), .ZN(n694) );
  XOR2_X1 U558 ( .A(KEYINPUT74), .B(n595), .Z(n514) );
  NOR2_X1 U559 ( .A1(n826), .A2(n825), .ZN(n515) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n693) );
  INV_X1 U561 ( .A(KEYINPUT89), .ZN(n700) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n717) );
  XNOR2_X1 U563 ( .A(n718), .B(n717), .ZN(n723) );
  OR2_X1 U564 ( .A1(G1384), .A2(n682), .ZN(n683) );
  XNOR2_X1 U565 ( .A(n687), .B(KEYINPUT64), .ZN(n692) );
  INV_X1 U566 ( .A(KEYINPUT94), .ZN(n763) );
  INV_X1 U567 ( .A(G2105), .ZN(n520) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n520), .ZN(n889) );
  BUF_X1 U569 ( .A(n685), .Z(G160) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U571 ( .A1(n891), .A2(G113), .ZN(n518) );
  AND2_X1 U572 ( .A1(n520), .A2(G2104), .ZN(n553) );
  NAND2_X1 U573 ( .A1(G101), .A2(n553), .ZN(n516) );
  XOR2_X1 U574 ( .A(n516), .B(KEYINPUT23), .Z(n517) );
  NAND2_X1 U575 ( .A1(n518), .A2(n517), .ZN(n524) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n519), .Z(n885) );
  NAND2_X1 U578 ( .A1(G137), .A2(n885), .ZN(n522) );
  NAND2_X1 U579 ( .A1(G125), .A2(n889), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n685) );
  XNOR2_X1 U582 ( .A(G2446), .B(G2443), .ZN(n534) );
  XOR2_X1 U583 ( .A(G2430), .B(KEYINPUT99), .Z(n526) );
  XNOR2_X1 U584 ( .A(G2454), .B(G2435), .ZN(n525) );
  XNOR2_X1 U585 ( .A(n526), .B(n525), .ZN(n530) );
  XOR2_X1 U586 ( .A(G2438), .B(G2427), .Z(n528) );
  XNOR2_X1 U587 ( .A(G1341), .B(G1348), .ZN(n527) );
  XNOR2_X1 U588 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U589 ( .A(n530), .B(n529), .Z(n532) );
  XNOR2_X1 U590 ( .A(KEYINPUT98), .B(G2451), .ZN(n531) );
  XNOR2_X1 U591 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U592 ( .A(n534), .B(n533), .ZN(n535) );
  AND2_X1 U593 ( .A1(n535), .A2(G14), .ZN(G401) );
  NAND2_X1 U594 ( .A1(G138), .A2(n885), .ZN(n540) );
  AND2_X1 U595 ( .A1(G102), .A2(n553), .ZN(n539) );
  NAND2_X1 U596 ( .A1(G114), .A2(n891), .ZN(n537) );
  NAND2_X1 U597 ( .A1(G126), .A2(n889), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n682) );
  AND2_X1 U600 ( .A1(n540), .A2(n682), .ZN(G164) );
  XOR2_X1 U601 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NOR2_X1 U602 ( .A1(G651), .A2(n632), .ZN(n642) );
  NAND2_X1 U603 ( .A1(G52), .A2(n642), .ZN(n544) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n542) );
  INV_X1 U605 ( .A(G651), .ZN(n545) );
  NOR2_X1 U606 ( .A1(G543), .A2(n545), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n650) );
  NAND2_X1 U608 ( .A1(G64), .A2(n650), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n551) );
  NOR2_X1 U610 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U611 ( .A1(G90), .A2(n646), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n632), .A2(n545), .ZN(n643) );
  NAND2_X1 U613 ( .A1(G77), .A2(n643), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n548), .Z(n549) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n549), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U619 ( .A1(G123), .A2(n889), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT18), .B(n552), .Z(n558) );
  NAND2_X1 U621 ( .A1(G99), .A2(n553), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G111), .A2(n891), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT77), .B(n556), .Z(n557) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n885), .A2(G135), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n920) );
  XNOR2_X1 U628 ( .A(G2096), .B(n920), .ZN(n561) );
  OR2_X1 U629 ( .A1(G2100), .A2(n561), .ZN(G156) );
  INV_X1 U630 ( .A(G57), .ZN(G237) );
  INV_X1 U631 ( .A(G132), .ZN(G219) );
  NAND2_X1 U632 ( .A1(G88), .A2(n646), .ZN(n563) );
  NAND2_X1 U633 ( .A1(G75), .A2(n643), .ZN(n562) );
  NAND2_X1 U634 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G50), .A2(n642), .ZN(n565) );
  NAND2_X1 U636 ( .A1(G62), .A2(n650), .ZN(n564) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U638 ( .A1(n567), .A2(n566), .ZN(G166) );
  NAND2_X1 U639 ( .A1(n646), .A2(G89), .ZN(n568) );
  XNOR2_X1 U640 ( .A(n568), .B(KEYINPUT4), .ZN(n570) );
  NAND2_X1 U641 ( .A1(G76), .A2(n643), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U643 ( .A(KEYINPUT5), .B(n571), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n650), .A2(G63), .ZN(n572) );
  XOR2_X1 U645 ( .A(KEYINPUT75), .B(n572), .Z(n574) );
  NAND2_X1 U646 ( .A1(n642), .A2(G51), .ZN(n573) );
  NAND2_X1 U647 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U648 ( .A(KEYINPUT6), .B(n575), .Z(n576) );
  NAND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U650 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT72), .ZN(n580) );
  XNOR2_X1 U654 ( .A(KEYINPUT10), .B(n580), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n835) );
  NAND2_X1 U656 ( .A1(n835), .A2(G567), .ZN(n581) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  NAND2_X1 U658 ( .A1(n646), .A2(G81), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n582), .B(KEYINPUT12), .ZN(n584) );
  NAND2_X1 U660 ( .A1(G68), .A2(n643), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT13), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G43), .A2(n642), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n650), .A2(G56), .ZN(n588) );
  XOR2_X1 U666 ( .A(KEYINPUT14), .B(n588), .Z(n589) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U668 ( .A(KEYINPUT73), .B(n591), .ZN(n1000) );
  INV_X1 U669 ( .A(n1000), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(G860), .ZN(G153) );
  INV_X1 U671 ( .A(G171), .ZN(G301) );
  NAND2_X1 U672 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G79), .A2(n643), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G54), .A2(n642), .ZN(n594) );
  NAND2_X1 U675 ( .A1(G92), .A2(n646), .ZN(n593) );
  NAND2_X1 U676 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n650), .A2(G66), .ZN(n595) );
  NOR2_X1 U678 ( .A1(n596), .A2(n514), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT15), .ZN(n993) );
  INV_X1 U681 ( .A(n993), .ZN(n614) );
  INV_X1 U682 ( .A(G868), .ZN(n661) );
  NAND2_X1 U683 ( .A1(n614), .A2(n661), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G91), .A2(n646), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G53), .A2(n642), .ZN(n603) );
  NAND2_X1 U687 ( .A1(G65), .A2(n650), .ZN(n602) );
  NAND2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U689 ( .A1(G78), .A2(n643), .ZN(n604) );
  XNOR2_X1 U690 ( .A(KEYINPUT69), .B(n604), .ZN(n605) );
  NOR2_X1 U691 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(KEYINPUT70), .ZN(G299) );
  NOR2_X1 U694 ( .A1(G286), .A2(n661), .ZN(n611) );
  NOR2_X1 U695 ( .A1(G299), .A2(G868), .ZN(n610) );
  NOR2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U697 ( .A(KEYINPUT76), .B(n612), .ZN(G297) );
  INV_X1 U698 ( .A(G559), .ZN(n616) );
  NOR2_X1 U699 ( .A1(G860), .A2(n616), .ZN(n613) );
  NOR2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U701 ( .A(KEYINPUT16), .B(n615), .Z(G148) );
  NAND2_X1 U702 ( .A1(n616), .A2(n993), .ZN(n617) );
  NAND2_X1 U703 ( .A1(n617), .A2(G868), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n1000), .A2(n661), .ZN(n618) );
  NAND2_X1 U705 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U706 ( .A1(G55), .A2(n642), .ZN(n621) );
  NAND2_X1 U707 ( .A1(G93), .A2(n646), .ZN(n620) );
  NAND2_X1 U708 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n643), .A2(G80), .ZN(n622) );
  XOR2_X1 U710 ( .A(KEYINPUT78), .B(n622), .Z(n623) );
  NOR2_X1 U711 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n650), .A2(G67), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(n660) );
  NAND2_X1 U714 ( .A1(G559), .A2(n993), .ZN(n627) );
  XNOR2_X1 U715 ( .A(n627), .B(n1000), .ZN(n658) );
  NOR2_X1 U716 ( .A1(G860), .A2(n658), .ZN(n628) );
  XOR2_X1 U717 ( .A(n660), .B(n628), .Z(G145) );
  NAND2_X1 U718 ( .A1(G49), .A2(n642), .ZN(n630) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U720 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U721 ( .A1(n650), .A2(n631), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U723 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G48), .A2(n642), .ZN(n636) );
  NAND2_X1 U725 ( .A1(G86), .A2(n646), .ZN(n635) );
  NAND2_X1 U726 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U727 ( .A1(n643), .A2(G73), .ZN(n637) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n637), .Z(n638) );
  NOR2_X1 U729 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n650), .A2(G61), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U732 ( .A1(G47), .A2(n642), .ZN(n645) );
  NAND2_X1 U733 ( .A1(G72), .A2(n643), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n646), .A2(G85), .ZN(n647) );
  XOR2_X1 U736 ( .A(KEYINPUT66), .B(n647), .Z(n648) );
  NOR2_X1 U737 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n650), .A2(G60), .ZN(n651) );
  NAND2_X1 U739 ( .A1(n652), .A2(n651), .ZN(G290) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(G288), .ZN(n657) );
  XNOR2_X1 U741 ( .A(G299), .B(G305), .ZN(n653) );
  XNOR2_X1 U742 ( .A(n653), .B(n660), .ZN(n654) );
  XNOR2_X1 U743 ( .A(G166), .B(n654), .ZN(n655) );
  XNOR2_X1 U744 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U745 ( .A(n657), .B(n656), .ZN(n908) );
  XNOR2_X1 U746 ( .A(n658), .B(n908), .ZN(n659) );
  NAND2_X1 U747 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G219), .A2(G220), .ZN(n668) );
  XNOR2_X1 U758 ( .A(KEYINPUT22), .B(n668), .ZN(n669) );
  NAND2_X1 U759 ( .A1(n669), .A2(G96), .ZN(n670) );
  NOR2_X1 U760 ( .A1(n670), .A2(G218), .ZN(n671) );
  XNOR2_X1 U761 ( .A(n671), .B(KEYINPUT79), .ZN(n841) );
  NAND2_X1 U762 ( .A1(n841), .A2(G2106), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G120), .A2(G69), .ZN(n672) );
  NOR2_X1 U764 ( .A1(G237), .A2(n672), .ZN(n673) );
  XNOR2_X1 U765 ( .A(KEYINPUT80), .B(n673), .ZN(n674) );
  NAND2_X1 U766 ( .A1(n674), .A2(G108), .ZN(n675) );
  XOR2_X1 U767 ( .A(KEYINPUT81), .B(n675), .Z(n840) );
  NAND2_X1 U768 ( .A1(G567), .A2(n840), .ZN(n676) );
  XNOR2_X1 U769 ( .A(KEYINPUT82), .B(n676), .ZN(n677) );
  NAND2_X1 U770 ( .A1(n678), .A2(n677), .ZN(n842) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U772 ( .A1(n842), .A2(n679), .ZN(n839) );
  NAND2_X1 U773 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  INV_X1 U775 ( .A(KEYINPUT65), .ZN(n761) );
  INV_X1 U776 ( .A(G1384), .ZN(n680) );
  AND2_X1 U777 ( .A1(G138), .A2(n680), .ZN(n681) );
  NAND2_X1 U778 ( .A1(n885), .A2(n681), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n684), .A2(n683), .ZN(n783) );
  NAND2_X1 U780 ( .A1(n685), .A2(G40), .ZN(n782) );
  INV_X1 U781 ( .A(n782), .ZN(n686) );
  NAND2_X1 U782 ( .A1(n783), .A2(n686), .ZN(n687) );
  XNOR2_X1 U783 ( .A(KEYINPUT86), .B(n692), .ZN(n705) );
  INV_X1 U784 ( .A(n705), .ZN(n719) );
  NAND2_X1 U785 ( .A1(n719), .A2(G2067), .ZN(n689) );
  BUF_X2 U786 ( .A(n692), .Z(n732) );
  NAND2_X1 U787 ( .A1(n732), .A2(G1348), .ZN(n688) );
  NAND2_X1 U788 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U789 ( .A(n690), .B(KEYINPUT88), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n732), .A2(G1341), .ZN(n696) );
  INV_X1 U791 ( .A(G1996), .ZN(n691) );
  XNOR2_X1 U792 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n1000), .A2(n697), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n702), .A2(n993), .ZN(n698) );
  NAND2_X1 U796 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n701), .B(n700), .ZN(n704) );
  OR2_X1 U798 ( .A1(n993), .A2(n702), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n711) );
  NAND2_X1 U800 ( .A1(G1956), .A2(n705), .ZN(n706) );
  XNOR2_X1 U801 ( .A(KEYINPUT87), .B(n706), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n719), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U803 ( .A(KEYINPUT27), .B(n707), .ZN(n708) );
  NOR2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n713) );
  INV_X1 U805 ( .A(G299), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U809 ( .A(n714), .B(KEYINPUT28), .Z(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U812 ( .A1(n719), .A2(n944), .ZN(n721) );
  INV_X1 U813 ( .A(G1961), .ZN(n966) );
  NAND2_X1 U814 ( .A1(n732), .A2(n966), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n727), .A2(G171), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n746) );
  NOR2_X1 U818 ( .A1(n732), .A2(G2084), .ZN(n750) );
  NOR2_X1 U819 ( .A1(n750), .A2(n747), .ZN(n724) );
  NAND2_X1 U820 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U822 ( .A1(G168), .A2(n726), .ZN(n729) );
  NOR2_X1 U823 ( .A1(G171), .A2(n727), .ZN(n728) );
  NOR2_X2 U824 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U825 ( .A(KEYINPUT31), .B(n730), .Z(n745) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n826), .ZN(n731) );
  XOR2_X1 U827 ( .A(KEYINPUT91), .B(n731), .Z(n734) );
  NOR2_X1 U828 ( .A1(n732), .A2(G2090), .ZN(n733) );
  NOR2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U830 ( .A1(n735), .A2(G303), .ZN(n737) );
  AND2_X1 U831 ( .A1(n745), .A2(n737), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n746), .A2(n736), .ZN(n740) );
  INV_X1 U833 ( .A(n737), .ZN(n738) );
  OR2_X1 U834 ( .A1(n738), .A2(G286), .ZN(n739) );
  AND2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U836 ( .A(n741), .B(KEYINPUT92), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n742), .A2(G8), .ZN(n744) );
  XOR2_X1 U838 ( .A(KEYINPUT32), .B(KEYINPUT93), .Z(n743) );
  XNOR2_X1 U839 ( .A(n744), .B(n743), .ZN(n819) );
  AND2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n749), .B(KEYINPUT90), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n750), .A2(G8), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n818) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  AND2_X1 U846 ( .A1(n818), .A2(n1001), .ZN(n753) );
  NAND2_X1 U847 ( .A1(n819), .A2(n753), .ZN(n758) );
  INV_X1 U848 ( .A(n1001), .ZN(n756) );
  NOR2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U851 ( .A1(n1003), .A2(n754), .ZN(n755) );
  OR2_X1 U852 ( .A1(n756), .A2(n755), .ZN(n757) );
  AND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U854 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U855 ( .A(n764), .B(n763), .ZN(n817) );
  NAND2_X1 U856 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U857 ( .A1(n826), .A2(n765), .ZN(n766) );
  XNOR2_X1 U858 ( .A(n766), .B(KEYINPUT95), .ZN(n815) );
  XNOR2_X1 U859 ( .A(G1981), .B(G305), .ZN(n991) );
  NAND2_X1 U860 ( .A1(G117), .A2(n891), .ZN(n768) );
  NAND2_X1 U861 ( .A1(G141), .A2(n885), .ZN(n767) );
  NAND2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n553), .A2(G105), .ZN(n769) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n769), .Z(n770) );
  NOR2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n889), .A2(G129), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n901) );
  NOR2_X1 U868 ( .A1(G1996), .A2(n901), .ZN(n918) );
  NAND2_X1 U869 ( .A1(G95), .A2(n553), .ZN(n775) );
  NAND2_X1 U870 ( .A1(G131), .A2(n885), .ZN(n774) );
  NAND2_X1 U871 ( .A1(n775), .A2(n774), .ZN(n779) );
  NAND2_X1 U872 ( .A1(G107), .A2(n891), .ZN(n777) );
  NAND2_X1 U873 ( .A1(G119), .A2(n889), .ZN(n776) );
  NAND2_X1 U874 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n881) );
  INV_X1 U876 ( .A(G1991), .ZN(n952) );
  NOR2_X1 U877 ( .A1(n881), .A2(n952), .ZN(n781) );
  AND2_X1 U878 ( .A1(G1996), .A2(n901), .ZN(n780) );
  NOR2_X1 U879 ( .A1(n781), .A2(n780), .ZN(n929) );
  NOR2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U881 ( .A(KEYINPUT83), .B(n784), .Z(n806) );
  XNOR2_X1 U882 ( .A(KEYINPUT85), .B(n806), .ZN(n785) );
  NOR2_X1 U883 ( .A1(n929), .A2(n785), .ZN(n809) );
  NOR2_X1 U884 ( .A1(G1986), .A2(G290), .ZN(n787) );
  AND2_X1 U885 ( .A1(n952), .A2(n881), .ZN(n786) );
  XNOR2_X1 U886 ( .A(KEYINPUT96), .B(n786), .ZN(n931) );
  NOR2_X1 U887 ( .A1(n787), .A2(n931), .ZN(n788) );
  XOR2_X1 U888 ( .A(KEYINPUT97), .B(n788), .Z(n789) );
  NOR2_X1 U889 ( .A1(n809), .A2(n789), .ZN(n790) );
  NOR2_X1 U890 ( .A1(n918), .A2(n790), .ZN(n791) );
  XNOR2_X1 U891 ( .A(n791), .B(KEYINPUT39), .ZN(n802) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n553), .A2(G104), .ZN(n792) );
  XNOR2_X1 U894 ( .A(n792), .B(KEYINPUT84), .ZN(n794) );
  NAND2_X1 U895 ( .A1(G140), .A2(n885), .ZN(n793) );
  NAND2_X1 U896 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n795), .ZN(n800) );
  NAND2_X1 U898 ( .A1(G116), .A2(n891), .ZN(n797) );
  NAND2_X1 U899 ( .A1(G128), .A2(n889), .ZN(n796) );
  NAND2_X1 U900 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n798), .Z(n799) );
  NOR2_X1 U902 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n801), .ZN(n902) );
  NOR2_X1 U904 ( .A1(n803), .A2(n902), .ZN(n935) );
  NAND2_X1 U905 ( .A1(n806), .A2(n935), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n802), .A2(n808), .ZN(n804) );
  NAND2_X1 U907 ( .A1(n803), .A2(n902), .ZN(n936) );
  NAND2_X1 U908 ( .A1(n804), .A2(n936), .ZN(n805) );
  NAND2_X1 U909 ( .A1(n805), .A2(n806), .ZN(n828) );
  INV_X1 U910 ( .A(n828), .ZN(n813) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n997) );
  NAND2_X1 U912 ( .A1(n997), .A2(n806), .ZN(n807) );
  AND2_X1 U913 ( .A1(n808), .A2(n807), .ZN(n811) );
  INV_X1 U914 ( .A(n809), .ZN(n810) );
  AND2_X1 U915 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U916 ( .A1(n813), .A2(n812), .ZN(n831) );
  NOR2_X1 U917 ( .A1(n991), .A2(n831), .ZN(n814) );
  AND2_X1 U918 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U919 ( .A1(n817), .A2(n816), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n819), .A2(n818), .ZN(n822) );
  NOR2_X1 U921 ( .A1(G2090), .A2(G303), .ZN(n820) );
  NAND2_X1 U922 ( .A1(G8), .A2(n820), .ZN(n821) );
  NAND2_X1 U923 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U924 ( .A1(n823), .A2(n826), .ZN(n827) );
  NOR2_X1 U925 ( .A1(G1981), .A2(G305), .ZN(n824) );
  XOR2_X1 U926 ( .A(n824), .B(KEYINPUT24), .Z(n825) );
  NOR2_X1 U927 ( .A1(n827), .A2(n515), .ZN(n829) );
  AND2_X1 U928 ( .A1(n829), .A2(n828), .ZN(n830) );
  OR2_X1 U929 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U930 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U932 ( .A1(n835), .A2(G2106), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n836), .B(KEYINPUT100), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U935 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U938 ( .A(G120), .B(KEYINPUT101), .ZN(G236) );
  XOR2_X1 U939 ( .A(G69), .B(KEYINPUT102), .Z(G235) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G325) );
  XNOR2_X1 U941 ( .A(KEYINPUT103), .B(G325), .ZN(G261) );
  XNOR2_X1 U942 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(n842), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U953 ( .A(G2084), .B(G2078), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1991), .B(G1976), .Z(n852) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1971), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n852), .B(n851), .ZN(n862) );
  XOR2_X1 U958 ( .A(G2474), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U959 ( .A(G1961), .B(KEYINPUT106), .ZN(n853) );
  XNOR2_X1 U960 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U961 ( .A(G1986), .B(G1981), .Z(n856) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1956), .ZN(n855) );
  XNOR2_X1 U963 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U964 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U965 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n859) );
  XNOR2_X1 U966 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U967 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G100), .A2(n553), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G112), .A2(n891), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U971 ( .A(n865), .B(KEYINPUT107), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G136), .A2(n885), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n889), .A2(G124), .ZN(n868) );
  XOR2_X1 U975 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  NOR2_X1 U976 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G103), .A2(n553), .ZN(n872) );
  NAND2_X1 U978 ( .A1(G139), .A2(n885), .ZN(n871) );
  NAND2_X1 U979 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G115), .A2(n891), .ZN(n874) );
  NAND2_X1 U981 ( .A1(G127), .A2(n889), .ZN(n873) );
  NAND2_X1 U982 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U984 ( .A1(n877), .A2(n876), .ZN(n922) );
  XOR2_X1 U985 ( .A(G162), .B(n922), .Z(n878) );
  XNOR2_X1 U986 ( .A(n920), .B(n878), .ZN(n900) );
  XOR2_X1 U987 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n880) );
  XNOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n879) );
  XNOR2_X1 U989 ( .A(n880), .B(n879), .ZN(n882) );
  XOR2_X1 U990 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U991 ( .A(G160), .B(G164), .ZN(n883) );
  XNOR2_X1 U992 ( .A(n884), .B(n883), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G106), .A2(n553), .ZN(n887) );
  NAND2_X1 U994 ( .A1(G142), .A2(n885), .ZN(n886) );
  NAND2_X1 U995 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U996 ( .A(KEYINPUT45), .B(n888), .Z(n896) );
  NAND2_X1 U997 ( .A1(n889), .A2(G130), .ZN(n890) );
  XNOR2_X1 U998 ( .A(n890), .B(KEYINPUT108), .ZN(n893) );
  NAND2_X1 U999 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U1000 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U1001 ( .A(n894), .B(KEYINPUT109), .Z(n895) );
  NOR2_X1 U1002 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U1003 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U1004 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n902), .B(n901), .Z(n903) );
  XNOR2_X1 U1006 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1008 ( .A(KEYINPUT112), .B(G286), .Z(n907) );
  XNOR2_X1 U1009 ( .A(G171), .B(n993), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(n907), .B(n906), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n1000), .B(n908), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(G401), .A2(n913), .ZN(n914) );
  AND2_X1 U1017 ( .A1(G319), .A2(n914), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n919), .Z(n933) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n921) );
  NAND2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1026 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1028 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1029 ( .A(KEYINPUT50), .B(n925), .Z(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  NAND2_X1 U1037 ( .A1(n939), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1038 ( .A(G2072), .B(G33), .Z(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT115), .B(n940), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G26), .B(G2067), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT116), .B(n943), .Z(n949) );
  XOR2_X1 U1043 ( .A(n944), .B(G27), .Z(n946) );
  XNOR2_X1 U1044 ( .A(G32), .B(G1996), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(KEYINPUT117), .B(n947), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(n950), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n951), .A2(G28), .ZN(n955) );
  XOR2_X1 U1050 ( .A(G25), .B(n952), .Z(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT114), .B(n953), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1053 ( .A(KEYINPUT53), .B(n956), .Z(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n957), .B(G34), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(G2084), .B(n958), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(G35), .B(G2090), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n963), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n964), .B(KEYINPUT55), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n965), .ZN(n1018) );
  XNOR2_X1 U1063 ( .A(n966), .B(G5), .ZN(n987) );
  XOR2_X1 U1064 ( .A(G1966), .B(G21), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G1986), .B(G24), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G22), .ZN(n967) );
  XNOR2_X1 U1067 ( .A(n967), .B(KEYINPUT124), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(G23), .B(G1976), .ZN(n968) );
  NOR2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1070 ( .A(KEYINPUT125), .B(n970), .ZN(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n973), .ZN(n974) );
  NAND2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n985) );
  XOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .Z(n976) );
  XNOR2_X1 U1075 ( .A(G4), .B(n976), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(G20), .B(G1956), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n980) );
  XNOR2_X1 U1079 ( .A(G6), .B(G1981), .ZN(n979) );
  NOR2_X1 U1080 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1081 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1082 ( .A(KEYINPUT60), .B(n983), .ZN(n984) );
  NOR2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(n988), .B(KEYINPUT61), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(n989), .ZN(n1019) );
  NOR2_X1 U1087 ( .A1(KEYINPUT123), .A2(n1019), .ZN(n1015) );
  XOR2_X1 U1088 ( .A(G168), .B(G1966), .Z(n990) );
  NOR2_X1 U1089 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1090 ( .A(KEYINPUT57), .B(n992), .Z(n999) );
  XNOR2_X1 U1091 ( .A(n993), .B(G1348), .ZN(n995) );
  XNOR2_X1 U1092 ( .A(G171), .B(G1961), .ZN(n994) );
  NAND2_X1 U1093 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1094 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1095 ( .A1(n999), .A2(n998), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(n1000), .B(G1341), .Z(n1011) );
  XNOR2_X1 U1097 ( .A(G299), .B(G1956), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G166), .B(G1971), .ZN(n1002) );
  NAND2_X1 U1099 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1100 ( .A(KEYINPUT120), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1101 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1102 ( .A(KEYINPUT121), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1103 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1104 ( .A(KEYINPUT122), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1105 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(KEYINPUT56), .A2(n1021), .ZN(n1014) );
  NOR2_X1 U1108 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1016), .ZN(n1017) );
  NOR2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1027) );
  INV_X1 U1111 ( .A(n1019), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(KEYINPUT123), .A2(n1020), .ZN(n1024) );
  INV_X1 U1113 ( .A(n1021), .ZN(n1022) );
  NAND2_X1 U1114 ( .A1(KEYINPUT56), .A2(n1022), .ZN(n1023) );
  NAND2_X1 U1115 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1116 ( .A1(n1025), .A2(G16), .ZN(n1026) );
  AND2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

